--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   10:46:38 07/09/2022
-- Design Name:   
-- Module Name:   E:/VHDL/Project/FinalProject/VM.TLB.Cache.Memory.Simulator/MainMemoryTest.vhd
-- Project Name:  VM.TLB.Cache.Memory.Simulator
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mainMemory
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MainMemoryTest IS
END MainMemoryTest;
 
ARCHITECTURE behavior OF MainMemoryTest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mainMemory
    PORT(
         outputData : OUT  std_logic_vector(31 downto 0);
         outputData2 : OUT  std_logic_vector(31 downto 0);
         PPN : OUT  std_logic_vector(3 downto 0);
         physicalAddressInput : IN  std_logic_vector(10 downto 0);
         virtualAddress : IN  std_logic_vector(15 downto 0);
         clock : IN  std_logic;
         controller : IN  std_logic;
         cache_type : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal physicalAddressInput : std_logic_vector(10 downto 0) := (others => '0');
   signal virtualAddress : std_logic_vector(15 downto 0) := (others => '0');
   signal clock : std_logic := '0';
   signal controller : std_logic := '0';
   signal cache_type : std_logic := '0';

 	--Outputs
   signal outputData : std_logic_vector(31 downto 0);
   signal outputData2 : std_logic_vector(31 downto 0);
   signal PPN : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clock_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: mainMemory PORT MAP (
          outputData => outputData,
          outputData2 => outputData2,
          PPN => PPN,
          physicalAddressInput => physicalAddressInput,
          virtualAddress => virtualAddress,
          clock => clock,
          controller => controller,
          cache_type => cache_type
        );

   -- Clock process definitions
   clock_process :process
   begin
		clock <= '0';
		wait for clock_period/2;
		clock <= '1';
		wait for clock_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clock_period*10;
		
      -- insert stimulus here 
		physicalAddressInput<="UUUUUUUUUUU";
		virtualAddress <="1111111011011111";
		controller <='1';
		cache_type <='U';
      wait;
   end process;

END;
