----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;



entity HardDisk is
    Port ( --PhysicalAddressIn : in  STD_LOGIC_VECTOR (10 downto 0);
           VirtualAddress : in  STD_LOGIC_VECTOR (15 downto 0);
           PhysicalAddressOut : out  STD_LOGIC_VECTOR (10 downto 0);
           outputData : out  STD_LOGIC_VECTOR (63 downto 0);
				cache_type : in std_logic; -- 0 --> direct , 1 --> 2 way
			  --controller : in std_logic; -- page table --> 0 
													-- datamemory --> 1 
				clock : in std_logic);
end HardDisk;

architecture Behavioral of HardDisk is
	type VirtualAdressInput is array (0 to 999) of std_logic_vector (15 downto 0);
	type PhysicalAdress is array (0 to 999) of std_logic_vector (10 downto 0);
	type DataTypeOutput is array (0 to 999) of std_logic_vector (31 downto 0);
	signal PAdress : PhysicalAdress := (0 => "10110111111", 1 => "00101111101", 2 => "01011001100",3 => "11101110100", 4 => "11100110110"
																	,5 => "10011001101",6 => "10000010110", 7 => "01100011110", 8 => "11101111011", 9 => "10010111000",10 => "00111111111",
																	11 => "01011001111", 12 => "01111111101",13 => "11101100111",14 => "00011000100",15 => "10100101101",16 => "10000111101",
																	17 => "10000000111",18 => "00011101000",19 => "00010011110", 20 => "01101101111",21 => "10001001111",22 => "10010101010", 23 => "11100100110"
																	,24 => "00110001100", 25 => "11000011111", 26 => "11010011010", 27 => "00000111010", 28 => "10011111100", 29 => "10011100101", 30 => "01111111101", 31 => "11100000001"
																	,32 => "10111101001",33 => "10110001111",34 => "10110001000",35 => "10101100110",36 => "10110110110",37 => "01111100111",38 => "10001101110"
																	,39 => "10100111111",40 => "10000011101",41 => "10001110111" ,42 => "00110000010",43 => "00100100010",44 =>"10110001010", 45 =>"10101110101",46 =>"11101000010"
																	,47 => "11000011100", 48 => "10100001000", 49 => "01111110010", 50 => "00100111000", 51 => "11011101111", 52 =>"01100110010",53 => "00111111100"
																	,54 => "10010001110",55 => "11111111011",56 => "10010100010",57 => "00011010010", 58 => "00011000110", 59 => "11010001010", 60 => "01101110000"
																	,61 => "01100000111", 62 => "00111000101", 63 => "11011011100", 64 => "11110101101", 65 => "11110111010", 66 => "10010101111", 67 => "01101000111"
																	,68 => "00010011100",69 => "11110011010", 70 => "00001111110", 71 => "11001010111", 72 => "00111110100", 73 => "01001111101", 74 => "11101000000"
																	,75 => "00010101011",76 => "00001111010", 77 => "00011100000", 78 => "10000000110", 79 => "01011111000", 80 => "11001110011", 81 => "00000010110"
																	,82 => "11010000000",83 => "00100101100", 84 => "10000111001", 85 => "00100001001", 86 => "01011001010", 87 => "01110111111", 88 => "01100111001"
																	,89 => "11010111100", 90 => "00100011000", 91 => "11110011011", 92 => "11101001100", 93 => "01011100001", 94 => "01111000100", 95 =>"00000001000"
																	,96 => "01101101110", 97 => "01000000001", 98 => "00000000111",99 => "01111100001",100 => "10000001110", 101 => "10111101101", 102 => "00000010011"
																	,103 => "10101101111",104 => "10010011100",105 => "00101111101",106 => "10011010101", 107 => "11101111010", 108 => "01111101111", 109 => "00011010010",
																	110 => "01000110000",111 => "11010110101", 112 => "00001001110",113 => "11101110000", 114 => "11110001000", 115 => "10010011001", 116 =>"10111010010",
																	117 => "01010010110", 118 => "10111000011", 119 => "01010001100", 120 => "11100010001", 121 => "10110111010", 122 => "01101101101", 123 => "11111110111", 124 => "11010110101", 125 => "00101110100", 126 => "01011111110", 127 => "10010100010", 128 => "00011000010", 129 => "10000100100", 130 => "11000000101", 131 => "10000111101"
																	,132 => "10000001010", 133 => "01100101000", 134 => "01111110111", 135 => "10100010101", 136 => "11111101100", 137 => "00000010100", 138 => "00010101000", 139 => "00000101010", 140 => "00011110111", 141 => "11011011000", 142 => "11011001101", 143 => "01101101100"
																	,144 => "00000001000", 145 => "11011101111", 146 => "11100110100", 147 => "10101001011", 148 => "11111100000", 149 => "00101010000", 150 =>"10101110110", 151 => "10010011111", 152 =>"00110110100", 153 => "10001110110", 154 => "01000111011", 155 => "10110111011", 156 => "10100001010", 157 => "01101010110", 158 => "00011110010", 159 => "11111100011"
																	,160 => "01010011101",161 => "10111011000", 162 => "00110010001", 163 => "11110110010", 164 => "10000000010", 165 => "00100010100", 166 => "01110100100", 167 => "01111111000", 168 => "00101000001", 169 => "10001010110", 170 => "01110011010", 171 => "11011100001", 172 => "01100011110", 173 => "01101101011", 174 => "11111001110", 175 => "11110100001", 176 => "10000010011", 177 => "00111010110", 178 => "01011111101", 179 => "11101101111", 180 => "00101001000", 181 => "01111001110"
																	,182 => "01001010111", 183 => "00101000000", 184 => "11011011011", 185 => "10101111001", 186 => "01001000011", 187 => "01000011110", 188 => "10111010110", 189 => "01010100111", 190 => "00010111110", 191 => "11100100011", 192 => "10101011000", 193 => "00010010111"
																	,194 => "11011110010", 195 => "10111001001", 196 => "10001011000", 197 => "00001111111", 198 => "10011001011", 199 => "11010001000", 200 => "11000101111", 201 => "01110110001", 202 => "11100010111", 203 => "10011101001", 204 => "10010101100", 205 =>"11111001100", 206 => "01110111000", 207 => "00010110100", 208 =>"00010110111", 209 => "11111000111", 210 => "01110000111", 211 => "01000101011", 212 => "00100000000", 213 => "01110101101", 214 => "00001011011", 215 => "01101101000", 216 => "01010100010"
																	,217 => "01100100000", 218 => "00010001100", 219 => "01000011010", 220 => "11011101011", 221 => "11000000011", 222 => "00110000111", 223 => "00001111001", 224 => "00010111000", 225 => "00000011100", 226 => "01011001110", 227 => "10111010101"
																	, 228 => "11010110111", 229 =>"01101001011", 230 => "11111101110", 231 => "00010000100", 232 => "01110010001", 233 => "00100000111", 234 => "11011000001", 235 => "01010010011", 236 => "11100010100", 237 => "00110010001", 238 => "01000110011", 239 => "10110101011"
																	, 240 => "11000001001", 241 => "00100110100", 242 => "10000001001", 243 => "11110101111", 244 => "11000101000", 245 => "01100011100", 246 => "00000100101", 247 => "10000110001", 248 => "10000001010", 249 => "11100101001", 250 => "11000000000", 251 => "00010011100"
																	, 252 => "00000110001", 253 => "10100010001", 254 => "10001110111", 255 => "11011101101", 256 =>"01111111111", 257 => "10011100101", 258 =>"11111001011", 259 =>"11101111101", 260 =>"00000101011", 261 => "11001010010", 262 => "01111111010", 263 =>"00010011110", 264 =>"01000111011", 265 => "01101010000"
																	,266 => "01110010001", 267 => "10101001111", 268 => "01111011101", 269 => "01010001111", 270 =>"00110101100", 271 => "11001001101", 272 =>"00011101010", 273 => "11110000001", 274 => "11101110000", 275 => "00001001000", 276 => "10110111000", 277 =>"10011010011", 278 =>"01111011010"
																	, 279 =>"10001000110", 280 => "11001110010", 281 =>"11000001000", 282 =>"00111110101", 283 =>"00001100100", 284 => "01010011000", 285 => "00100111111", 286 => "11011001110", 287 => "11000111000", 288 => "01001001111", 289 => "01100100001", 290 => "01011010011", 291 => "01101010111", 292 => "10000111011", 293 => "10100010010", 294 => "10000010001", 295 => "11111010101", 296 => "00100111011"
																	,297 => "11011010101", 298 => "01100110100", 299 => "00110010011", 
																	300 => "11000101111", 301 => "01110110001", 302 => "11100010111", 303 => "10011101001", 304 => "10010101100", 305 =>"11111001100", 306 => "01110111000", 307 => "00010110100", 308 => "00010110111", 309 => "11111000111", 310 => "01110000111",311 => "01000101011", 312 => "00100000000", 313 => "01110101101", 314 => "00001011011", 315 => "01101101000", 316 => "01010100010"
																	,317 => "01100100000", 318 => "00010001100", 319 => "01000011010", 320 => "11011101011", 321 => "11000000011", 322 => "00110000111", 323 => "00001111001", 324 => "00010111000", 325 => "00000011100", 326 => "01011001110", 327 => "10111010101"
																	, 328 => "11010110111", 329 =>"01101001011", 330 => "11111101110", 331 => "00010000100", 332 => "01110010001", 333 => "00100000111", 334 => "11011000001", 335 => "01010010011", 336 => "11100010100", 337 => "00110010001", 338 => "01000110011", 339 => "10110101011"
																	, 340 => "11000001001", 341 => "00100110100", 342 => "10000001001", 343 => "11110101111", 344 => "11000101000", 345 => "01100011100", 346 => "00000100101", 347 => "10000110001", 348 => "10000001010", 349 => "11100101001", 350 => "11000000000", 351 => "00010011100"
																	, 352 => "00000110001", 353 => "10100010001", 354 => "10001110111", 355 => "11011101101", 356 =>"01111111111", 357 => "10011100101", 358 =>"11111001011", 359 =>"11101111101", 360 =>"00000101011", 361 => "11001010010", 362 => "01111111010", 363 =>"00010011110", 364 =>"01000111011", 365 => "01101010000"
																	,366 => "01110010001", 367 => "10101001111", 368 => "01111011101", 369 => "01010001111", 370 =>"00110101100", 371 => "11001001101", 372 =>"00011101010", 373 => "11110000001", 374 => "11101110000", 375 => "00001001000", 376 => "10110111000", 377 =>"10011010011", 378 =>"01111011010"
																	,379 =>"10001000110", 380 => "11001110010", 381 =>"11000001000", 382 =>"00111110101", 383 =>"00001100100", 384 => "01010011000", 385 => "00100111111", 386 => "11011001110", 387 => "11000111000", 388 => "01001001111", 389 => "01100100001", 390 => "01011010011", 391 => "01101010111", 392 => "10000111011", 393 => "10100010010", 394 => "10000010001", 395 => "11111010101", 396 => "00100111011"
																	,397 => "11011010101", 398 => "01100110100", 399 => "00110010011",
																	400 => "11000101111", 401 => "01110110001", 402 => "11100010111", 403 => "10011101001", 404 => "10010101100", 405 =>"11111001100", 406 => "01110111000", 407 => "00010110100", 408 => "00010110111", 409 => "11111000111", 410 => "01110000111",411 => "01000101011", 412 => "00100000000", 413 => "01110101101", 414 => "00001011011", 415 => "01101101000", 416 => "01010100010"
																	,417 => "01100100000", 418 => "00010001100", 419 => "01000011010", 420 => "11011101011", 421 => "11000000011", 422 => "00110000111", 423 => "00001111001", 424 => "00010111000", 425 => "00000011100", 426 => "01011001110", 427 => "10111010101"
																	, 428 => "11010110111", 429 =>"01101001011", 430 => "11111101110", 431 => "00010000100", 432 => "01110010001", 433 => "00100000111", 434 => "11011000001", 435 => "01010010011", 436 => "11100010100", 437 => "00110010001", 438 => "01000110011", 439 => "10110101011"
																	, 440 => "11000001001", 441 => "00100110100", 442 => "10000001001", 443 => "11110101111", 444 => "11000101000", 445 => "01100011100", 446 => "00000100101", 447 => "10000110001", 448 => "10000001010", 449 => "11100101001", 450 => "11000000000", 451 => "00010011100"
																	, 452 => "00000110001", 453 => "10100010001", 454 => "10001110111", 455 => "11011101101", 456 =>"01111111111", 457 => "10011100101", 458 =>"11111001011", 459 =>"11101111101", 460 =>"00000101011", 461 => "11001010010", 462 => "01111111010", 463 =>"00010011110", 464 =>"01000111011", 465 => "01101010000"
																	,466 => "01110010001", 467 => "10101001111", 468 => "01111011101", 469 => "01010001111", 470 =>"00110101100", 471 => "11001001101", 472 =>"00011101010", 473 => "11110000001", 474 => "11101110000", 475 => "00001001000", 476 => "10110111000", 477 =>"10011010011", 478 =>"01111011010"
																	,479 =>"10001000110", 480 => "11001110010", 481 =>"11000001000", 482 =>"00111110101", 483 =>"00001100100", 484 => "01010011000", 485 => "00100111111", 486 => "11011001110", 487 => "11000111000", 488 => "01001001111", 489 => "01100100001", 490 => "01011010011", 491 => "01101010111", 492 => "10000111011", 493 => "10100010010", 494 => "10000010001", 495 => "11111010101", 496 => "00100111011"
																	,497 => "11011010101", 498 => "01100110100", 499 => "00110010011",
																	500 => "11000101111", 501 => "01110110001", 502 => "11100010111", 503 => "10011101001", 504 => "10010101100", 505 =>"11111001100", 506 => "01110111000", 507 => "00010110100", 508 => "00010110111", 509 => "11111000111", 510 => "01110000111", 511 => "01000101011", 512 => "00100000000", 513 => "01110101101", 514 => "00001011011", 515 => "01101101000", 516 => "01010100010"
																	,517 => "01100100000", 518 => "00010001100", 519 => "01000011010", 520 => "11011101011", 521 => "11000000011", 522 => "00110000111", 523 => "00001111001", 524 => "00010111000", 525 => "00000011100", 526 => "01011001110", 527 => "10111010101"
																	, 528 => "11010110111", 529 =>"01101001011", 530 => "11111101110", 531 => "00010000100", 532 => "01110010001", 533 => "00100000111", 534 => "11011000001", 535 => "01010010011", 536 => "11100010100", 537 => "00110010001", 538 => "01000110011", 539 => "10110101011"
																	, 540 => "11000001001", 541 => "00100110100", 542 => "10000001001", 543 => "11110101111", 544 => "11000101000", 545 => "01100011100", 546 => "00000100101", 547 => "10000110001", 548 => "10000001010", 549 => "11100101001", 550 => "11000000000", 551 => "00010011100"
																	, 552 => "00000110001", 553 => "10100010001", 554 => "10001110111", 555 => "11011101101", 556 =>"01111111111", 557 => "10011100101", 558 =>"11111001011", 559 =>"11101111101", 560 =>"00000101011", 561 => "11001010010", 562 => "01111111010", 563 =>"00010011110", 564 =>"01000111011", 565 => "01101010000"
																	,566 => "01110010001", 567 => "10101001111", 568 => "01111011101", 569 => "01010001111", 570 =>"00110101100", 571 => "11001001101", 572 =>"00011101010", 573 => "11110000001", 574 => "11101110000", 575 => "00001001000", 576 => "10110111000", 577 =>"10011010011", 578 =>"01111011010"
																	,579 =>"10001000110", 580 => "11001110010", 581 =>"11000001000", 582 =>"00111110101", 583 =>"00001100100", 584 => "01010011000", 585 => "00100111111", 586 => "11011001110", 587 => "11000111000", 588 => "01001001111", 589 => "01100100001", 590 => "01011010011", 591 => "01101010111", 592 => "10000111011", 593 => "10100010010", 594 => "10000010001", 595 => "11111010101", 596 => "00100111011"
																	,597 => "11011010101", 598 => "01100110100", 599 => "00110010011",			
																	600 => "11000101111", 601 => "01110110001", 602 => "11100010111", 603 => "10011101001", 604 => "10010101100", 605 =>"11111001100", 606 => "01110111000", 607 => "00010110100", 608 => "00010110111", 609 => "11111000111", 610 => "01110000111",611 => "01000101011", 612 => "00100000000", 613 => "01110101101", 614 => "00001011011", 615 => "01101101000", 616 => "01010100010"
																	,617 => "01100100000", 618 => "00010001100", 619 => "01000011010", 620 => "11011101011", 621 => "11000000011", 622 => "00110000111", 623 => "00001111001", 624 => "00010111000", 625 => "00000011100", 626 => "01011001110", 627 => "10111010101"
																	, 628 => "11010110111", 629 =>"01101001011", 630 => "11111101110", 631 => "00010000100", 632 => "01110010001", 633 => "00100000111", 634 => "11011000001", 635 => "01010010011", 636 => "11100010100", 637 => "00110010001", 638 => "01000110011", 639 => "10110101011"
																	, 640 => "11000001001", 641 => "00100110100", 642 => "10000001001", 643 => "11110101111", 644 => "11000101000", 645 => "01100011100", 646 => "00000100101", 647 => "10000110001", 648 => "10000001010", 649 => "11100101001", 650 => "11000000000", 651 => "00010011100"
																	, 652 => "00000110001", 653 => "10100010001", 654 => "10001110111", 655 => "11011101101", 656 =>"01111111111", 657 => "10011100101", 658 =>"11111001011", 659 =>"11101111101", 660 =>"00000101011", 661 => "11001010010", 662 => "01111111010", 663 =>"00010011110", 664 =>"01000111011", 665 => "01101010000"
																	,666 => "01110010001", 667 => "10101001111", 668 => "01111011101", 669 => "01010001111", 670 =>"00110101100", 671 => "11001001101", 672 =>"00011101010", 673 => "11110000001", 674 => "11101110000", 675 => "00001001000", 676 => "10110111000", 677 =>"10011010011", 678 =>"01111011010"
																	,679 =>"10001000110", 680 => "11001110010", 681 =>"11000001000", 682 =>"00111110101", 683 =>"00001100100", 684 => "01010011000", 685 => "00100111111", 686 => "11011001110", 687 => "11000111000", 688 => "01001001111", 689 => "01100100001", 690 => "01011010011", 691 => "01101010111", 692 => "10000111011", 693 => "10100010010", 694 => "10000010001", 695 => "11111010101", 696 => "00100111011"
																	,697 => "11011010101", 698 => "01100110100", 699 => "00110010011",
																	700 => "11000101111", 701 => "01110110001", 702 => "11100010111", 703 => "10011101001", 704 => "10010101100", 705 =>"11111001100", 706 => "01110111000", 707 => "00010110100", 708 => "00010110111", 709 => "11111000111", 710 => "01110000111",711 => "01000101011", 712 => "00100000000", 713 => "01110101101", 714 => "00001011011", 715 => "01101101000", 716 => "01010100010"
																	,717 => "01100100000", 718 => "00010001100", 719 => "01000011010", 720 => "11011101011", 721 => "11000000011", 722 => "00110000111", 723 => "00001111001", 724 => "00010111000", 725 => "00000011100", 726 => "01011001110", 727 => "10111010101"
																	, 728 => "11010110111", 729 =>"01101001011", 730 => "11111101110", 731 => "00010000100", 732 => "01110010001", 733 => "00100000111", 734 => "11011000001", 735 => "01010010011", 736 => "11100010100", 737 => "00110010001", 738 => "01000110011", 739 => "10110101011"
																	, 740 => "11000001001", 741 => "00100110100", 742 => "10000001001", 743 => "11110101111", 744 => "11000101000", 745 => "01100011100", 746 => "00000100101", 747 => "10000110001", 748 => "10000001010", 749 => "11100101001", 750 => "11000000000", 751 => "00010011100"
																	, 752 => "00000110001", 753 => "10100010001", 754 => "10001110111", 755 => "11011101101", 756 =>"01111111111", 757 => "10011100101", 758 =>"11111001011", 759 =>"11101111101", 760 =>"00000101011", 761 => "11001010010", 762 => "01111111010", 763 =>"00010011110", 764 =>"01000111011", 765 => "01101010000"
																	,766 => "01110010001", 767 => "10101001111", 768 => "01111011101", 769 => "01010001111", 770 =>"00110101100", 771 => "11001001101", 772 =>"00011101010", 773 => "11110000001", 774 => "11101110000", 775 => "00001001000", 776 => "10110111000", 777 =>"10011010011", 778 =>"01111011010"
																	,779 =>"10001000110", 780 => "11001110010", 781 =>"11000001000", 782 =>"00111110101", 783 =>"00001100100", 784 => "01010011000", 785 => "00100111111", 786 => "11011001110", 787 => "11000111000", 788 => "01001001111", 789 => "01100100001", 790 => "01011010011", 791 => "01101010111", 792 => "10000111011", 793 => "10100010010", 794 => "10000010001", 795 => "11111010101", 796 => "00100111011"
																	,797 => "11011010101", 798 => "01100110100", 799 => "00110010011",
																	800 => "11000101111", 801 => "01110110001", 802 => "11100010111", 803 => "10011101001", 804 => "10010101100", 805 =>"11111001100", 806 => "01110111000", 807 => "00010110100", 808 => "00010110111", 809 => "11111000111", 810 => "01110000111",811 => "01000101011", 812 => "00100000000", 813 => "01110101101", 814 => "00001011011", 815 => "01101101000", 816 => "01010100010"
																	,817 => "01100100000", 818 => "00010001100", 819 => "01000011010", 820 => "11011101011", 821 => "11000000011", 822 => "00110000111", 823 => "00001111001", 824 => "00010111000", 825 => "00000011100", 826 => "01011001110", 827 => "10111010101"
																	, 828 => "11010110111", 829 =>"01101001011", 830 => "11111101110", 831 => "00010000100", 832 => "01110010001", 833 => "00100000111", 834 => "11011000001", 835 => "01010010011", 836 => "11100010100", 837 => "00110010001", 838 => "01000110011", 839 => "10110101011"
																	, 840 => "11000001001", 841 => "00100110100", 842 => "10000001001", 843 => "11110101111", 844 => "11000101000", 845 => "01100011100", 846 => "00000100101", 847 => "10000110001", 848 => "10000001010", 849 => "11100101001", 850 => "11000000000", 851 => "00010011100"
																	, 852 => "00000110001", 853 => "10100010001", 854 => "10001110111", 855 => "11011101101", 856 =>"01111111111", 857 => "10011100101", 858 =>"11111001011", 859 =>"11101111101", 860 =>"00000101011", 861 => "11001010010", 862 => "01111111010", 863 =>"00010011110", 864 =>"01000111011", 865 => "01101010000"
																	,866 => "01110010001", 867 => "10101001111", 868 => "01111011101", 869 => "01010001111", 870 =>"00110101100", 871 => "11001001101", 872 =>"00011101010", 873 => "11110000001", 874 => "11101110000", 875 => "00001001000", 876 => "10110111000", 877 =>"10011010011", 878 =>"01111011010"
																	,879 =>"10001000110", 880 => "11001110010", 881 =>"11000001000", 882 =>"00111110101", 883 =>"00001100100", 884 => "01010011000", 885 => "00100111111", 886 => "11011001110", 887 => "11000111000", 888 => "01001001111", 889 => "01100100001", 890 => "01011010011", 891 => "01101010111", 892 => "10000111011", 893 => "10100010010", 894 => "10000010001", 895 => "11111010101", 896 => "00100111011"
																	,897 => "11011010101", 898 => "01100110100", 899 => "00110010011",
																	900 => "11000101111", 901 => "01110110001", 902 => "11100010111", 903 => "10011101001", 904 => "10010101100", 905 =>"11111001100", 906 => "01110111000", 907 => "00010110100", 908 => "00010110111", 909 => "11111000111", 910 => "01110000111",911 => "01000101011", 912 => "00100000000", 913 => "01110101101", 914 => "00001011011", 915 => "01101101000", 916 => "01010100010"
																	,917 => "01100100000", 918 => "00010001100", 919 => "01000011010", 920 => "11011101011", 921 => "11000000011", 922 => "00110000111", 923 => "00001111001", 924 => "00010111000", 925 => "00000011100", 926 => "01011001110", 927 => "10111010101"
																	, 928 => "11010110111", 929 =>"01101001011", 930 => "11111101110", 931 => "00010000100", 932 => "01110010001", 933 => "00100000111", 934 => "11011000001", 935 => "01010010011", 936 => "11100010100", 937 => "00110010001", 938 => "01000110011", 939 => "10110101011"
																	, 940 => "11000001001", 941 => "00100110100", 942 => "10000001001", 943 => "11110101111", 944 => "11000101000", 945 => "01100011100", 946 => "00000100101", 947 => "10000110001", 948 => "10000001010", 949 => "11100101001", 950 => "11000000000", 951 => "00010011100"
																	, 952 => "00000110001", 953 => "10100010001", 954 => "10001110111", 955 => "11011101101", 956 =>"01111111111", 957 => "10011100101", 958 =>"11111001011", 959 =>"11101111101", 960 =>"00000101011", 961 => "11001010010", 962 => "01111111010", 963 =>"00010011110", 964 =>"01000111011", 965 => "01101010000"
																	,966 => "01110010001", 967 => "10101001111", 968 => "01111011101", 969 => "01010001111", 970 =>"00110101100", 971 => "11001001101", 972 =>"00011101010", 973 => "11110000001", 974 => "11101110000", 975 => "00001001000", 976 => "10110111000", 977 =>"10011010011", 978 =>"01111011010"
																	,979 =>"10001000110", 980 => "11001110010", 981 =>"11000001000", 982 =>"00111110101", 983 =>"00001100100", 984 => "01010011000", 985 => "00100111111", 986 => "11011001110", 987 => "11000111000", 988 => "01001001111", 989 => "01100100001", 990 => "01011010011", 991 => "01101010111", 992 => "10000111011", 993 => "10100010010", 994 => "10000010001", 995 => "11111010101", 996 => "00100111011"
																	,997 => "11011010101", 998 => "01100110100", 999 => "00110010011");
	
	
	signal VAdress : VirtualAdressInput := (0 => "1111111010111111", 1 => "1111110011111101", 2 => "1111110101001100",3 => "1111111111110100", 4 => "1111111110110110"
																	,5 => "1111100110011111",6 => "1000001011111110", 7 => "0110011111101110", 8 => "1110111111111011", 9 => "1001011100111110",10 => "1111110011111111",
																	11 => "1111100110011111", 12 => "1111000111111101",13 => "1111001111100111",14 => "1111000001000100",15 => "1111001010101101",16 => "1111001000011101",
																	17 => "1111100000001111",18 => "1111000011101000",19 => "1111000000011110", 20 => "1111000101101111",21 => "1111001001001111",22 => "1111001001011010", 23 => "1111001110010011"
																	,24 => "1111001100011001", 25 => "0000011000011111", 26 => "0000011010011010", 27 => "0000000000111010", 28 => "0000010011111100", 29 => "0000000011100101", 30 => "0000000111111101", 31 => "0000011100000001"
																   ,32 => "1111101111010011",33 => "1011011111100111",34 => "1011001111101000",35 => "1010110110111111",36 => "1011111110110110",37 => "0111110111110111",38 => "1011111100110110"
																	,39 => "1111101001111111",40 => "1001111110001101",41 => "1011111001110111" ,42 => "0011011111100010",43 => "0010010111111001",44 =>"1011001111101010", 45 =>"1010111011111101",46 =>"1110100111110010"
																	,47 => "1111110000111001", 48 => "1010111111001000", 49 => "0111110111111010", 50 => "0101111110111000", 51 => "1101110111111111", 52 =>"0110110111111010",53 => "0011111111111100"
																	,54 => "1111110010001101",55 => "1111111111111011",56 => "1011111101010010",57 => "0001111111010010", 58 => "0001111111100010", 59 => "1111111010001010", 60 => "1111110111110000"
																	,61 => "1111101100001111", 62 => "0011100111110101", 63 => "1101101110011111", 64 => "1111010111111110", 65 => "1111011111111010", 66 => "1111111010101111", 67 => "0110111111100111"
																	,68 => "1111100010011100",69 => "1111001111111010", 70 => "0011111100111110", 71 => "1100101100111011", 72 => "0011111001110100", 73 => "1001111001111101", 74 => "1110000011001100"
																	,75 => "0011001101101011",76 => "0000111101111010", 77 => "0001110011100000", 78 => "1000000011100110", 79 => "0101111100111000", 80 => "1100111100111011", 81 => "1101100000010110"
																	,82 => "1101000010011000",83 => "0010110110101100", 84 => "1000011100111001", 85 => "0010011001100001", 86 => "0101101001101010", 87 => "0111101111001111", 88 => "0110111100111001"
																	,89 => "1101011100111100", 90 => "0010011100111000", 91 => "1111001110011011", 92 => "1110100111011100", 93 => "0101110011100001", 94 => "0111100110010100", 95 =>"0011001100001000"
																	,96 => "0110110110011110", 97 => "0100100110000001", 98 => "0000100110000111",99 => "0111110011100001",																	
																	100 => "1000000110011110", 101 => "1011110011110110", 102 => "0011001100010011"
																	,103 => "1010110111001111",104 => "1001001110011100",105 => "0010111110011101",106 => "1001110011010101", 107 => "1110111001111010", 108 => "0111101110011111", 109 => "0001101010011010",
																	110 => "0100011001010100",111 => "1101010101010101", 112 => "0001001110101010",113 => "1101010110111000", 114 => "1101010110001000", 115 => "1001001110101001", 116 =>"1011010101010010",
																	117 => "0101001011011111", 118 => "1011100001111111", 119 => "0101000110011111", 120 => "1110101010010001", 121 => "1010101011011010", 122 => "1010100110101101", 123 => "1110101011110111", 124 => "1101010101010101", 125 => "0010110101010100", 126 => "0101110101011110", 127 => "1001010011010010", 128 => "0010101001100010", 129 => "1000101100100100", 130 => "1100001010100101", 131 => "1001010100011101"
																	,132 => "1001010100001010", 133 => "0110100100101000", 134 => "0111010111110111", 135 => "1010011010010101", 136 => "1010011111101100", 137 => "0010110000010100", 138 => "0101010010101000", 139 => "0010110000101010", 140 => "0001111011010101", 141 => "1101101101010100", 142 =>"1101101010100101", 143 => "0110110101010100"
																	,144 => "0000101010001000", 145 => "1101110101010111", 146 => "1101010100110100", 147 => "1010101011001011", 148 => "1010101111100000", 149 => "0010101001001000", 150 =>"1010110101011110", 151 => "1001001101010111", 152 =>"0011011001010100", 153 => "1000110101010110", 154 => "0100101010011011", 155 => "1011011010101011", 156 => "1010101010001010", 157 => "1010100101010110", 158 => "0010101001110010", 159 => "1110101011100011"
																	,160 => "0101001110011111",161 => "1011101010101000", 162 => "0011010101010001", 163 => "1101010110110010", 164 => "1010101000000010", 165 => "0010010101000100", 166 => "0111010101010100", 167 => "0111101010111000", 168 => "0010100010101001", 169 => "1001010110101010", 170 => "0110011010101010", 171 => "1101110010101001", 172 => "1010100110001110", 173 => "1010100101101011", 174 => "1110101011100110", 175 => "1110101011010001", 176 => "1000101010000011", 177 => "0101010011110110", 178 => "0101110101011101", 179 => "1110110111010111", 180 => "0010100101011000", 181 => "0111010101100110"
																	,182 => "0101010110101011", 183 => "0010100101010000", 184 => "1101101010101011", 185 => "1010111010101001", 186 => "1010100100100011", 187 => "0100011010101110", 188 => "1011010101010110", 189 => "0101010101010011", 190 => "0010111010101110", 191 => "1110010011010101", 192 => "1010101100101010", 193 => "0010011010100111"
																	,194 => "1101111001011111", 195 => "1011010101001001", 196 => "1010101001011000", 197 => "0000111010101111", 198 => "1010101001101011", 199 => "1101010101001000", 																	
																	200 => "1100010110101011", 201 => "0111010101011001", 202 => "1110101010010111", 203 => "1001101010101001", 204 => "1001010110101010", 205 =>"1110101011001100", 206 => "1010100111011000", 207 => "1010100010110100", 208 =>"0010101001010111", 209 => "1111010101000111", 210 => "0111010101000011", 211 => "0101010100101011", 212 => "0010000101010000", 213 => "0111010110101010", 214 => "0001011010101011", 215 => "0110101010110100", 216 => "0101010010101010"
																	,217 => "0110010010101000", 218 => "0010011011001100", 219 => "0101101100011010", 220 => "1101110110110101", 221 => "1100001101100011", 222 => "0011001101100111", 223 => "0001111011011001", 224 => "0001011101101000", 225 => "0001101100011100", 226 => "0101101101100110", 227 => "1011101101010101"
																	, 228 => "1101011011101111", 229 =>"0110100101110110", 230 => "1111101101101110", 231 => "1101100010000100", 232 => "0111011010010001", 233 => "1101100010000111", 234 => "1101101101100001", 235 => "1101100101010011", 236 => "1110010100110110", 237 => "1101100110010001", 238 => "0100011001110110", 239 => "1011010101110110"
																	, 240 => "1100000100111011", 241 => "1101100100110100", 242 => "1010110000001001", 243 => "1111010111101101", 244 => "1101101100101000", 245 => "0110001111011000", 246 => "0000100101110110", 247 => "1000011001110110", 248 => "1101101000001010", 249 => "1110101001110110", 250 => "1101101100000000", 251 => "1101100010011100"
																	, 252 => "0000011000111011", 253 => "1101101010001001", 254 => "1001110111101101", 255 => "1101110110110101", 256 =>"1101100111111111", 257 => "1101101001100101", 258 =>"1101101111001011", 259 =>"1101101110111101", 260 =>"1101100000101011", 261 => "1101101101010010", 262 => "1101100111111010", 263 =>"1101100001001110", 264 =>"1101100100111011", 265 => "1101100110101000"
																	,266 => "0111001000101111", 267 => "1101101010100111", 268 => "0111101101011101", 269 => "0101001101100111", 270 =>"1101100110101100", 271 => "1101101101001101", 272 =>"1101100011101010", 273 => "1101101111000001", 274 => "1101101101110000", 275 => "1101100001001000", 276 => "1101101011011000", 277 =>"1101101001101011", 278 =>"1101100111011010"
																	, 279 =>"1000100011011011", 280 => "1111011000110010", 281 =>"1100001011011000", 282 =>"0011101101110101", 283 =>"1101100001100100", 284 => "1101100101011000", 285 => "1101100010011111", 286 => "1101101101100110", 287 => "1101101000111000", 288 => "1101100001001111", 289 => "1101100110010001", 290 => "1101100101101011", 291 => "1101100110101011", 292 => "1000011101110110", 293 => "1010010010110110", 294 => "1000010001110110", 295 => "1111010101110110", 296 => "0010011101110110"
																	,297 => "1101101010111011", 298 => "0110011011011010", 299 => "0011011011010011", 																																		
																	300 => "0000011000101111", 301 => "0000001110110001", 302 => "1110001011100000", 303 => "0000010011101001", 304 => "0000001001010110", 305 =>"0000011111001100", 306 => "0111011100000000", 307 => "0000000010110100", 308 => "0001011010000011", 309 => "1111100010000011", 310 => "0110000010000111",311 => "0100010101000001", 312 => "0010000000000000", 313 => "0111010100000101", 314 => "0001010000001011", 315 => "0110100000101000", 316 => "0101010000000010"
																	,317 => "0000001100100000", 318 => "0000000010001100", 319 => "0100001101000000", 320 => "0000011011101011", 321 => "1100000001100000", 322 => "0000000110000111", 323 => "0000111100100000", 324 => "0000000010111000", 325 => "0000001100000100", 326 => "0101100100000110", 327 => "1010000011010101"
																	, 328 => "0000011010110111", 329 =>"0000001101001011", 330 => "1111110111000000", 331 => "0000000010000100", 332 => "0000000111000001", 333 => "0000000100000111", 334 => "1101100000100000", 335 => "0101001001000001", 336 => "1100000100010100", 337 => "0010000010010001", 338 => "0100010000010011", 339 => "1010000010101011"
																	, 340 => "0000011000001001", 341 => "0000000100110100", 342 => "1000000100100000", 343 => "0000011110101111", 344 => "1100010100000000", 345 => "0000001100011100", 346 => "0000010010100000", 347 => "1000010000001001", 348 => "1000000000001010", 349 => "1000001100101001", 350 => "1000000100000000", 351 => "0001001000001100"
																	, 352 => "0000000000110001", 353 => "0000010100010001", 354 => "1000111011100000", 355 => "0000011011101101", 356 =>"0000000111111111", 357 => "0000000011100101", 358 =>"1111100101100000", 359 =>"1110111000001101", 360 =>"0000101010000001", 361 => "1000001001010010", 362 => "0111000001111010", 363 =>"0001001100000110", 364 =>"0100010000011011", 365 => "0110101000000000"
																	,366 => "0000001110010001", 367 => "0000010101001111", 368 => "0111101110100000", 369 => "0000001010001111", 370 =>"0011010110000000", 371 => "0000011001001101", 372 =>"0001110101000000", 373 => "1100000011000001", 374 => "1110100000110000", 375 => "0000100000001000", 376 => "1011011000001000", 377 =>"1001000001010011", 378 =>"0111000001011010"
																	,379 =>"0000010001000110", 380 => "0000011001110010", 381 =>"1100000100000000", 382 =>"0000000111110101", 383 =>"0000000000110100", 384 => "0000001010011000", 385 => "0010011111100000", 386 => "1101100110000010", 387 => "1100010000011000", 388 => "0100100110000011", 389 => "0100000100100001", 390 => "0101000001010011", 391 => "0110101011000001", 392 => "1000010000011011", 393 => "1010000000010010", 394 => "1000001000000001", 395 => "1110000011010101", 396 => "0010010000011011"
																	,397 => "0100110110101011", 398 => "0000011001101001", 399 => "0011001001100001",																	
																	400 => "1011111000101111", 401 => "1011101110110001", 402 => "1110001011110111", 403 => "1001110101111001", 404 => "1010111010101100", 405 =>"1111100101111100", 406 => "0111011110111000", 407 => "0001010111110100", 408 => "0001011011110111", 409 => "1101111111000111", 410 => "0111000101110111",411 => "0110111000101011", 412 => "0101110100000000", 413 => "0111010110111101", 414 => "0001011101011011", 415 => "0110101111101000", 416 => "0101010101110010"
																	,417 => "1011110110010000", 418 => "0101110010001100", 419 => "0100101110011010", 420 => "1101110111101011", 421 => "1101111000000011", 422 => "0011101110000111", 423 => "0010111001111001", 424 => "0001011110111000", 425 => "0000101110011100", 426 => "0101101011101110", 427 => "1011101111010101"
																	, 428 => "1011111010110111", 429 =>"0110110111001011", 430 => "1111110111101110", 431 => "0001010111000100", 432 => "1011101110010001", 433 => "0010010111000111", 434 => "1101101011100001", 435 => "0101010111010011", 436 => "1110101110010100", 437 => "0011010111010001", 438 => "0101011100110011", 439 => "1101110110101011"
																	, 440 => "1011111000001001", 441 => "0010101110110100", 442 => "1001011100001001", 443 => "1101111110101111", 444 => "1100010101111000", 445 => "0110010111011100", 446 => "0001011100100101", 447 => "1000101110110001", 448 => "1000101110001010", 449 => "1110101110101001", 450 => "1100000101110000", 451 => "0101110010011100"
																	, 452 => "1011100000110001", 453 => "1010010111010001", 454 => "1001011101110111", 455 => "1101111011101101", 456 =>"0111111011111111", 457 => "1001110010111111", 458 =>"1111101011101011", 459 =>"1110111101111101", 460 =>"0001011100101011", 461 => "1100101010111010", 462 => "0111111101111010", 463 =>"0010111010011110", 464 =>"0100011110111011", 465 => "0101111101010000"
																	,466 => "1011101110010001", 467 => "1010101011101111", 468 => "0111011111011101", 469 => "0101010111001111", 470 =>"0011011011101100", 471 => "1100101011101101", 472 =>"0010111011101010", 473 => "1111010111000001", 474 => "1110111011110000", 475 => "0010111001001000", 476 => "1010111110111000", 477 =>"1010111011010011", 478 =>"0111101110111010"
																	,479 =>"1011110001000110", 480 => "1100111011110010", 481 =>"1100010111001000", 482 =>"0011101111110101", 483 =>"0000110101110100", 484 => "0101010111011000", 485 => "0010011110111111", 486 => "1101101011101110", 487 => "1101011100111000", 488 => "0100101111001111", 489 => "0111011100100001", 490 => "0101111011010011", 491 => "0111011101010111", 492 => "1000010111111011", 493 => "1010010111010010", 494 => "1000101110010001", 495 => "1111101011110101", 496 => "0010010111111011"
																	,497 => "1011111011010101", 498 => "1011101100110100", 499 => "1011100110010011",																	
																	500 => "0011111000101111", 501 => "0111010011110001", 502 => "1110001001110111", 503 => "1001100111101001", 504 => "1001010100111100", 505 =>"1110011111001100", 506 => "0011101110111000", 507 => "0011100010110100", 508 => "0011100010110111", 509 => "1100111111000111", 510 => "0100111110000111", 511 => "0100001110101011", 512 => "0010001110000000", 513 => "0111000111101101", 514 => "0000111001011011", 515 => "0100111101101000", 516 => "0101010001110010"
																	,517 => "0011101100100000", 518 => "0001000111001100", 519 => "0100011100011010", 520 => "1101110011101011", 521 => "1100000011100011", 522 => "0000111110000111", 523 => "0011100001111001", 524 => "0011100010111000", 525 => "0011100000011100", 526 => "0001111011001110", 527 => "1001110111010101"
																	, 528 => "0011111010110111", 529 =>"0110001111001011", 530 => "1111100111101110", 531 => "0001001110000100", 532 => "0111001000011101", 533 => "0001110100000111", 534 => "0011111011000001", 535 => "0001111010010011", 536 => "0011111100010100", 537 => "0001110110010001", 538 => "0100111000110011", 539 => "1010011110101011"
																	, 540 => "0011111000001001", 541 => "0010011001110100", 542 => "1000000111001001", 543 => "1111000111101111", 544 => "1100010100001110", 545 => "0001111100011100", 546 => "0011100000100101", 547 => "0011110000110001", 548 => "0011110000001010", 549 => "0011111100101001", 550 => "1100111000000000", 551 => "0000011110011100"
																	, 552 => "0011100000110001", 553 => "1010000011110001", 554 => "1000001111110111", 555 => "1100011111101101", 556 =>"0111111001111111", 557 => "1001110011100101", 558 =>"0011111111001011", 559 =>"1100111101111101", 560 =>"0011100000101011", 561 => "1100111001010010", 562 => "0011101111111010", 563 =>"0000011110011110", 564 =>"0100001110111011", 565 => "0110001111010000"
																	,566 => "0011101110010001", 567 => "1010100110011111", 568 => "0111001111011101", 569 => "0101000111001111", 570 =>"0011010001111100", 571 => "1100111001001101", 572 =>"0011100011101010", 573 => "0011111110000001", 574 => "0011111101110000", 575 => "0011100001001000", 576 => "1001110110111000", 577 =>"1001101000111011", 578 =>"0100111111011010"
																	,579 =>"0011110001000110", 580 => "1100110011110010", 581 =>"1100000011101000", 582 =>"0011111000111101", 583 =>"0000110010000111", 584 => "0101001110011000", 585 => "0011100100111111", 586 => "1001111011001110", 587 => "0011111000111000", 588 => "0011101001001111", 589 => "0011101100100001", 590 => "0001111011010011", 591 => "0110011101010111", 592 => "1000000111111011", 593 => "1010000111010010", 594 => "1000011100010001", 595 => "1111100011110101", 596 => "0010011100111011"
																	,597 => "0011111011010101", 598 => "0110010011110100", 599 => "0011001001111111",																	
														      	600 => "0101111000101111", 601 => "0101101110110001", 602 => "0101111100010111", 603 => "0101110011101001", 604 => "0101110010101100", 605 =>"0101111111001100", 606 => "0101101110111000", 607 => "0101100010110100", 608 => "0101100010110111", 609 => "0101111111000111", 610 => "0101101110000111",611 => "0101101000101011", 612 => "0101100100000000", 613 => "0101101110101101", 614 => "0101100001011011", 615 => "0101101101101000", 616 => "0101101010100010"
																	,617 => "0101101100100000", 618 => "0101100010001100", 619 => "0101101000011010", 620 => "0101111011101011", 621 => "0101111000000011", 622 => "0101100110000111", 623 => "0101100001111001", 624 => "0101100010111000", 625 => "0101100000011100", 626 => "0101101011001110", 627 => "0101110111010101"
																	, 628 => "0101111010110111", 629 =>"0101101101001011", 630 => "0101111111101110", 631 => "0101100010000100", 632 => "0101101110010001", 633 => "0101100100000111", 634 => "0101111011000001", 635 => "0100101110010011", 636 => "0101111100010100", 637 => "0101100110010001", 638 => "0101101000110011", 639 => "0101110110101011"
																	, 640 => "0101111000001001", 641 => "0101100100110100", 642 => "0101110000001001", 643 => "0101111110101111", 644 => "0101111000101000", 645 => "0101101100011100", 646 => "0101100000100101", 647 => "1001011000110001", 648 => "0101110000001010", 649 => "0101111100101001", 650 => "0101111000000000", 651 => "0101100010011100"
																	, 652 => "0000011000111111", 653 => "0101110100010001", 654 => "0101110001110111", 655 => "0101111011101101", 656 =>"0101101111111111", 657 => "0101110011100101", 658 =>"0101111111001011", 659 =>"0101111101111101", 660 =>"0101100000101011", 661 => "0101111001010010", 662 => "0101101111111010", 663 =>"0101100010011110", 664 =>"0101101000111011", 665 => "0101101101010000"
																	,666 => "0101101110010001", 667 => "0101110101001111", 668 => "0101101111011101", 669 => "0101101010001111", 670 =>"0101100110101100", 671 => "0101111001001101", 672 =>"0101100011101010", 673 => "0101111110000001", 674 => "0101111101110000", 675 => "0101100001001000", 676 => "0101110110111000", 677 =>"0101110011010011", 678 =>"0101101111011010"
																	,679 =>"0101110001000110", 680 => "0101111001110010", 681 =>"1010111000001000", 682 =>"0101100111110101", 683 =>"0101100001100100", 684 => "0101101010011000", 685 => "0101100100111111", 686 => "0101111011001110", 687 => "0101111000111000", 688 => "0101101001001111", 689 => "0101101100100001", 690 => "0101101011010011", 691 => "0101101101010111", 692 => "0101110000111011", 693 => "0101110100010010", 694 => "0101110000010001", 695 => "0101111111010101", 696 => "0101100100111011"
																	,697 => "0101111011010101", 698 => "0101101100110100", 699 => "0101100110010011",																	
												    				700 => "1001011000101111", 701 => "1001001110110001", 702 => "1001011100010111", 703 => "1001010011101001", 704 => "1001010010101100", 705 =>"1001011111001100", 706 => "1001001110111000", 707 => "1001000010110100", 708 => "1001000010110111", 709 => "1001011111000111", 710 => "1001001110000111",711 => "1001001000101011", 712 => "1001000100000000", 713 => "1001001110101101", 714 => "1001000001011011", 715 => "1001001101101000", 716 => "1001001010100010"
																	,717 => "1001001100100000", 718 => "1001000010001100", 719 => "1001001000011010", 720 => "1001011011101011", 721 => "1001011000000011", 722 => "1001000110000111", 723 => "1001000001111001", 724 => "1001000010111000", 725 => "1001000000011100", 726 => "1001001011001110", 727 => "1001010111010101"
																	, 728 => "1001011010110111", 729 =>"1001001101001011", 730 => "1001011111101110", 731 => "1001000010000100", 732 => "1001001110010001", 733 => "1001000100000111", 734 => "1001011011000001", 735 => "1001001010010011", 736 => "1001011100010100", 737 => "1001000110010001", 738 => "1001001000110011", 739 => "1001010110101011"
																	, 740 => "1001011000001001", 741 => "1001000100110100", 742 => "1001010000001001", 743 => "1001011110101111", 744 => "1001011000101000", 745 => "1001001100011100", 746 => "1001000000100101", 747 => "1001010000110001", 748 => "1001010000001010", 749 => "1001011100101001", 750 => "1001011000000000", 751 => "1001000010011100"
																	, 752 => "1001000000110001", 753 => "1001010100010001", 754 => "1001010001110111", 755 => "1001011011101101", 756 =>"1001001111111111", 757 => "1001010011100101", 758 =>"1001011111001011", 759 =>"1001011101111101", 760 =>"1001000000101011", 761 => "1001011001010010", 762 => "1001001111111010", 763 =>"1001000010011110", 764 =>"1001001000111011", 765 => "1001001101010000"
																	,766 => "1001001110010001", 767 => "1001010101001111", 768 => "1001001111011101", 769 => "1001001010001111", 770 =>"1001000110101100", 771 => "1001011001001101", 772 =>"1001000011101010", 773 => "1001011110000001", 774 => "1001011101110000", 775 => "1001000001001000", 776 => "1001010110111000", 777 =>"1001010011010011", 778 =>"1001001111011010"
																	,779 =>"1001010001000110", 780 => "1001011001110010", 781 =>"1001011000001000", 782 =>"1001000111110101", 783 =>"1001000001100100", 784 => "1001001010011000", 785 => "1001000100111111", 786 => "1001011011001110", 787 => "1001011000111000", 788 => "1001001001001111", 789 => "1001001100100001", 790 => "1001001011010011", 791 => "1001001101010111", 792 => "1001010000111011", 793 => "1001010100010010", 794 => "1001010000010001", 795 => "1001011111010101", 796 => "1001000100111011"
																	,797 => "1001011011010101", 798 => "1001001100110100", 799 => "1001000110010011",																
																	800 => "1001011000101111", 801 => "1001001110110001", 802 => "1100101100010111", 803 => "1001010011101001", 804 => "1001010010101100", 805 =>"1001011111001100", 806 => "1001001110111000", 807 => "1001000010110100", 808 => "1001000010110111", 809 => "1001011111000111", 810 => "1001001110000111",811 => "1001001000101011", 812 => "1001000100000000", 813 => "1001001110101101", 814 => "1001000001011011", 815 => "1001001101101000", 816 => "1001001010100010"
																	,817 => "1001001100100000", 818 => "1001000010001100", 819 => "1001001000011010", 820 => "1001011011101011", 821 => "1001011000000011", 822 => "1001000110000111", 823 => "1001000001111001", 824 => "1001000010111000", 825 => "1001000000011100", 826 => "1001001011001110", 827 => "1001010111010101"
																	, 828 => "1001011010110111", 829 =>"1001001101001011", 830 => "1001011111101110", 831 => "1001000010000100", 832 => "1001001110010001", 833 => "1001000100000111", 834 => "1001011011000001", 835 => "1001001010010011", 836 => "1001011100010100", 837 => "1001000110010001", 838 => "1001001000110011", 839 => "1001010110101011"
																	, 840 => "1001011000001001", 841 => "1001000100110100", 842 => "1001010000001001", 843 => "1001011110101111", 844 => "1001011000101000", 845 => "1001001100011100", 846 => "1001000000100101", 847 => "1001010000110001", 848 => "1001010000001010", 849 => "1001011100101001", 850 => "1001011000000000", 851 => "1001000010011100"
																	, 852 => "1001000000110001", 853 => "1001010100010001", 854 => "1001010001110111", 855 => "1001011011101101", 856 =>"1001001111111111", 857 => "1001010011100101", 858 =>"1001011111001011", 859 =>"1001011101111101", 860 =>"1001000000101011", 861 => "1001011001010010", 862 => "1001001111111010", 863 =>"1001000010011110", 864 =>"1001001000111011", 865 => "1001001101010000"
																	,866 => "1001001110010001", 867 => "1001010101001111", 868 => "1001001111011101", 869 => "1001001010001111", 870 =>"1001000110101100", 871 => "1001011001001101", 872 =>"1001000011101010", 873 => "1001011110000001", 874 => "1001011101110000", 875 => "1001000001001000", 876 => "1001010110111000", 877 =>"1001010011010011", 878 =>"1001001111011010"
																	,879 =>"1001010001000110", 880 => "1001011001110010", 881 =>"1001011000001000", 882 =>"1001000111110101", 883 =>"1001000001100100", 884 => "1001001010011000", 885 => "1001000100111111", 886 => "1001011011001110", 887 => "1001011000111000", 888 => "1001001001001111", 889 => "1001001100100001", 890 => "1001001011010011", 891 => "1001001101010111", 892 => "1001010000111011", 893 => "1001010100010010", 894 => "1001010000010001", 895 => "1001011111010101", 896 => "1001000100111011"
																	,897 => "1001011011010101", 898 => "1001001100110100", 899 => "1001000110010011",
																	900 => "0000111000101111", 901 => "0111011000100001", 902 => "1110001011100001", 903 => "1001110100100001", 904 => "1001010110000001", 905 =>"0000111111001100", 906 => "0111011100000001", 907 => "0001011010000001", 908 => "0000100010110111", 909 => "1110000111000111", 910 => "0000101110000111",911 => "0000101000101011", 912 => "0000010100000000", 913 => "0000101110101101", 914 => "0000100001011011", 915 => "0000101101101000", 916 => "0000101010100010"
																	,917 => "0000101100100000", 918 => "0001000110000001", 919 => "0100001101000001", 920 => "1101110101100001", 921 => "1100000001100001", 922 => "0000100110000111", 923 => "0000111100100001", 924 => "0001011100000001", 925 => "0000100000011100", 926 => "0100001011001110", 927 => "1000010111010101"
																	, 928 => "0000111010110111", 929 =>"0110100101100001", 930 => "1111110111000001", 931 => "0001000010000001", 932 => "0111001000100001", 933 => "0000100100000111", 934 => "1101100000100001", 935 => "0101001001100001", 936 => "0000111100010100", 937 => "0000010110010001", 938 => "0000101000110011", 939 => "0000110110101011"
																	, 940 => "0000111000001001", 941 => "0010011010000001", 942 => "1000000100100001", 943 => "1111010111100001", 944 => "1100010100000001", 945 => "0000101100011100", 946 => "0000010010100001", 947 => "1000011000100001", 948 => "0000110000001010", 949 => "0000111100101001", 950 => "0000111000000000", 951 => "0000100010011100"
																	, 952 => "0000100000110001", 953 => "1010001000100001", 954 => "1000111011100001", 955 => "1101110110100001", 956 =>"0111111111100001", 957 => "0000110011100101", 958 =>"1111100101100001", 959 =>"1110111110100001", 960 =>"0000100000101011", 961 => "0000111001010010", 962 => "0000101111111010", 963 =>"0000100010011110", 964 =>"0100001000111011", 965 => "0000101101010000"
																	,966 => "0000101110010001", 967 => "1010100111100001", 968 => "0111101110100001", 969 => "0101000111100001", 970 =>"0011010110000001", 971 => "0000111001001101", 972 =>"0001110101000001", 973 => "1111000000100001", 974 => "0000111101110000", 975 => "0000100001001000", 976 => "0000110110111000", 977 =>"0000110011010011", 978 =>"0000011111011010"
																	,979 =>"0000110001000110", 980 => "1100111001000001", 981 =>"1100000100000001", 982 =>"0011111010100001", 983 =>"0000110010000001", 984 => "0000101010011000", 985 => "0010011111100001", 986 => "1101100111000001", 987 => "0000111000111000", 988 => "0000101001001111", 989 => "0000101100100001", 990 => "0000101011010011", 991 => "0000011101010111", 992 => "0000110000111011", 993 => "0000110100010010", 994 => "0000110000010001", 995 => "0000111111010101", 996 => "0000100100111011"
																	,997 => "0000111011010101", 998 => "0110011010000001", 999 => "0011001001100001");
	
	
	
	
	
	
	
	
	signal DataOutput1 : DataTypeOutput := (0 => "11111110110111111111111011011111", 1 => "11111100101111011111110010111101", 2 => "11111101011001101111110101100110",3 => "11111111101110101111111110111010", 4 => "11111111100110111111111110011011"
																	,5 => "11111001100111111111100110011111",6 => "10000010111111101000001011111110", 7 => "01100111111011100110011111101110", 8 => "11101111111110111110111111111011", 9 => "10010111001111101001011100111110",10 => "11111100111111111111110011111111",
																	11 => "11111001100111111111100110011111", 12 => "11110001111111011111000111111101",13 => "11110011111001111111001111100111",14 => "11110000010001001111000001000100",15 => "11110010101011011111001010101101",16 => "11110010000111011111001000011101",
																	17 => "11111000000011111111100000001111",18 => "11110000111010001111000011101000",19 => "11110000000111101111000000011110", 20 => "11110001011011111111000101101111",21 => "11110010010011111111001001001111",22 => "11110010010110101111001001011010", 23 => "11110011100100111111001110010011"
																	,24 => "11110011000110011111001100011001", 25 => "00000110000111110000011000011111", 26 => "00000110100110100000011010011010", 27 => "00000000001110100000000000111010", 28 => "00000100111111000000010011111100", 29 => "00000000111001010000000011100101", 30 => "00000001111111010000000111111101", 31 => "00000111000000010000011100000001"
																   ,32 => "11111011110100111111101111010011",33 => "10110111111001111011011111100111",34 => "10110011111010001011001111101000",35 => "10101101101111111010110110111111",36 => "10111111101101101011111110110110",37 => "01111101111101110111110111110111",38 => "10111111001101101011111100110110"
																	,39 => "11111010011111111111101001111111",40 => "10011111100011011001111110001101",41 => "10111110011101111011111001110111" ,42 => "00110111111000100011011111100010",43 => "00100101111110010010010111111001",44 =>"10110011111010101011001111101010", 45 =>"10101110111111011010111011111101",46 =>"11101001111100101110100111110010"
																	,47 => "11111100001110011111110000111001", 48 => "10101111110010001010111111001000", 49 => "01111101111110100111110111111010", 50 => "01011111101110000101111110111000", 51 => "11011101111111111101110111111111", 52 =>"01101101111110100110110111111010",53 => "00111111111111000011111111111100"
																	,54 => "11111100100011011111110010001101",55 => "11111111111110111111111111111011",56 => "10111111010100101011111101010010",57 => "00011111110100100001111111010010", 58 => "00011111111000100001111111100010", 59 => "11111110100010101111111010001010", 60 => "11111101111100001111110111110000"
																	,61 => "11111011000011111111101100001111", 62 => "00111001111101010011100111110101", 63 => "11011011100111111101101110011111", 64 => "11110101111111101111010111111110", 65 => "11110111111110101111011111111010", 66 => "11111110101011111111111010101111", 67 => "01101111111001110110111111100111"
																	,68 => "11111000100111001111100010011100",69 => "11110011111110101111001111111010", 70 => "00111111001111100011111100111110", 71 => "11001011001110111100101100111011", 72 => "00111110011101000011111001110100", 73 => "10011110011111011001111001111101", 74 => "11100000110011001110000011001100"
																	,75 => "00110011011010110011001101101011",76 => "00001111011110100000111101111010", 77 => "00011100111000000001110011100000", 78 => "10000000111001101000000011100110", 79 => "01011111001110000101111100111000", 80 => "11001111001110111100111100111011", 81 => "11011000000101101101100000010110"
																	,82 => "11010000100110001101000010011000",83 => "00101101101011000010110110101100", 84 => "10000111001110011000011100111001", 85 => "00100110011000010010011001100001", 86 => "01011010011010100101101001101010", 87 => "01111011110011110111101111001111", 88 => "01101111001110010110111100111001"
																	,89 => "11010111001111001101011100111100", 90 => "00100111001110000010011100111000", 91 => "11110011100110111111001110011011", 92 => "11101001110111001110100111011100", 93 => "01011100111000010101110011100001", 94 => "01111001100101000111100110010100", 95 =>"00110011000010000011001100001000"
																	,96 => "01101101100111100110110110011110", 97 => "01001001100000010100100110000001", 98 => "00001001100001110000100110000111",99 => "01111100111000010111110011100001",																	
																	100 => "10000001100111101000000110011110", 101 => "10111100111101101011110011110110", 102 => "00110011000100110011001100010011"
																	,103 => "10101101110011111010110111001111",104 => "10010011100111001001001110011100",105 => "00101111100111010010111110011101",106 => "10011100110101011001110011010101", 107 => "11101110011110101110111001111010", 108 => "01111011100111110111101110011111", 109 => "00011010100110100001101010011010",
																	110 => "01000110010101000100011001010100",111 => "11010101010101011101010101010101", 112 => "00010011101010100001001110101010",113 => "11010101101110001101010110111000", 114 => "11010101100010001101010110001000", 115 => "10010011101010011001001110101001", 116 =>"10110101010100101011010101010010",
																	117 => "01010010110111110101001011011111", 118 => "10111000011111111011100001111111", 119 => "01010001100111110101000110011111", 120 => "11101010100100011110101010010001", 121 => "10101010110110101010101011011010", 122 => "10101001101011011010100110101101", 123 => "11101010111101111110101011110111", 124 => "11010101010101011101010101010101", 125 => "00101101010101000010110101010100", 126 => "01011101010111100101110101011110", 127 => "10010100110100101001010011010010", 128 => "00101010011000100010101001100010", 129 => "10001011001001001000101100100100", 130 => "11000010101001011100001010100101", 131 => "10010101000111011001010100011101"
																	,132 => "10010101000010101001010100001010", 133 => "01101001001010000110100100101000", 134 => "01110101111101110111010111110111", 135 => "10100110100101011010011010010101", 136 => "10100111111011001010011111101100", 137 => "00101100000101000010110000010100", 138 => "01010100101010000101010010101000", 139 => "00101100001010100010110000101010", 140 => "00011110110101010001111011010101", 141 => "11011011010101001101101101010100", 142 =>"11011010101001011101101010100101", 143 => "01101101010101000110110101010100"
																	,144 => "00001010100010000000101010001000", 145 => "11011101010101111101110101010111", 146 => "11010101001101001101010100110100", 147 => "10101010110010111010101011001011", 148 => "10101011111000001010101111100000", 149 => "00101010010010000010101001001000", 150 =>"10101101010111101010110101011110", 151 => "10010011010101111001001101010111", 152 =>"00110110010101000011011001010100", 153 => "10001101010101101000110101010110", 154 => "01001010100110110100101010011011", 155 => "10110110101010111011011010101011", 156 => "10101010100010101010101010001010", 157 => "10101001010101101010100101010110", 158 => "00101010011100100010101001110010", 159 => "11101010111000111110101011100011"
																	,160 => "01010011100111110101001110011111",161 => "10111010101010001011101010101000", 162 => "00110101010100010011010101010001", 163 => "11010101101100101101010110110010", 164 => "10101010000000101010101000000010", 165 => "00100101010001000010010101000100", 166 => "01110101010101000111010101010100", 167 => "01111010101110000111101010111000", 168 => "00101000101010010010100010101001", 169 => "10010101101010101001010110101010", 170 => "01100110101010100110011010101010", 171 => "11011100101010011101110010101001", 172 => "10101001100011101010100110001110", 173 => "10101001011010111010100101101011", 174 => "11101010111001101110101011100110", 175 => "11101010110100011110101011010001", 176 => "10001010100000111000101010000011", 177 => "01010100111101100101010011110110", 178 => "01011101010111010101110101011101", 179 => "11101101110101111110110111010111", 180 => "00101001010110000010100101011000", 181 => "01110101011001100111010101100110"
																	,182 => "01010101101010110101010110101011", 183 => "00101001010100000010100101010000", 184 => "11011010101010111101101010101011", 185 => "10101110101010011010111010101001", 186 => "10101001001000111010100100100011", 187 => "01000110101011100100011010101110", 188 => "10110101010101101011010101010110", 189 => "01010101010100110101010101010011", 190 => "00101110101011100010111010101110", 191 => "11100100110101011110010011010101", 192 => "10101011001010101010101100101010", 193 => "00100110101001110010011010100111"
																	,194 => "11011110010111111101111001011111", 195 => "10110101010010011011010101001001", 196 => "10101010010110001010101001011000", 197 => "00001110101011110000111010101111", 198 => "10101010011010111010101001101011", 199 => "11010101010010001101010101001000", 																	
																	200 => "11000101101010111100010110101011", 201 => "01110101010110010111010101011001", 202 => "11101010100101111110101010010111", 203 => "10011010101010011001101010101001", 204 => "10010101101010101001010110101010", 205 =>"11101010110011001110101011001100", 206 => "10101001110110001010100111011000", 207 => "10101000101101001010100010110100", 208 =>"00101010010101110010101001010111", 209 => "11110101010001111111010101000111", 210 => "01110101010000110111010101000011", 211 => "01010101001010110101010100101011", 212 => "00100001010100000010000101010000", 213 => "01110101101010100111010110101010", 214 => "00010110101010110001011010101011", 215 => "01101010101101000110101010110100", 216 => "01010100101010100101010010101010"
																	,217 => "01100100101010000110010010101000", 218 => "00100110110011000010011011001100", 219 => "01011011000110100101101100011010", 220 => "11011101101101011101110110110101", 221 => "11000011011000111100001101100011", 222 => "00110011011001110011001101100111", 223 => "00011110110110010001111011011001", 224 => "00010111011010000001011101101000", 225 => "00011011000111000001101100011100", 226 => "01011011011001100101101101100110", 227 => "10111011010101011011101101010101"
																	,228 => "11010110111011111101011011101111", 229 =>"01101001011101100110100101110110", 230 => "11111011011011101111101101101110", 231 => "11011000100001001101100010000100", 232 => "01110110100100010111011010010001", 233 => "11011000100001111101100010000111", 234 => "11011011011000011101101101100001", 235 => "11011001010100111101100101010011", 236 => "11100101001101101110010100110110", 237 => "11011001100100011101100110010001", 238 => "01000110011101100100011001110110", 239 => "10110101011101101011010101110110"
																	,240 => "11000001001110111100000100111011", 241 => "11011001001101001101100100110100", 242 => "10101100000010011010110000001001", 243 => "11110101111011011111010111101101", 244 => "11011011001010001101101100101000", 245 => "01100011110110000110001111011000", 246 => "00001001011101100000100101110110", 247 => "10000110011101101000011001110110", 248 => "11011010000010101101101000001010", 249 => "11101010011101101110101001110110", 250 => "11011011000000001101101100000000", 251 => "11011000100111001101100010011100"
																	,252 => "00000110001110110000011000111011", 253 => "11011010100010011101101010001001", 254 => "10011101111011011001110111101101", 255 => "11011101101101011101110110110101", 256 =>"11011001111111111101100111111111", 257 => "11011010011001011101101001100101", 258 =>"11011011110010111101101111001011", 259 =>"11011011101111011101101110111101", 260 =>"11011000001010111101100000101011", 261 => "11011011010100101101101101010010", 262 => "11011001111110101101100111111010", 263 =>"11011000010011101101100001001110", 264 =>"11011001001110111101100100111011", 265 => "11011001101010001101100110101000"
																	,266 => "01110010001011110111001000101111", 267 => "11011010101001111101101010100111", 268 => "01111011010111010111101101011101", 269 => "01010011011001110101001101100111", 270 =>"11011001101011001101100110101100", 271 => "11011011010011011101101101001101", 272 =>"11011000111010101101100011101010", 273 => "11011011110000011101101111000001", 274 => "11011011011100001101101101110000", 275 => "11011000010010001101100001001000", 276 => "11011010110110001101101011011000", 277 =>"11011010011010111101101001101011", 278 =>"11011001110110101101100111011010"
																	,279 =>"10001000110110111000100011011011", 280 => "11110110001100101111011000110010", 281 =>"11000010110110001100001011011000", 282 =>"00111011011101010011101101110101", 283 =>"11011000011001001101100001100100", 284 => "11011001010110001101100101011000", 285 => "11011000100111111101100010011111", 286 => "11011011011001101101101101100110", 287 => "11011010001110001101101000111000", 288 => "11011000010011111101100001001111", 289 => "11011001100100011101100110010001", 290 => "11011001011010111101100101101011", 291 => "11011001101010111101100110101011", 292 => "10000111011101101000011101110110", 293 => "10100100101101101010010010110110", 294 => "10000100011101101000010001110110", 295 => "11110101011101101111010101110110", 296 => "00100111011101100010011101110110"
																	,297 => "11011010101110111101101010111011", 298 => "01100110110110100110011011011010", 299 => "00110110110100110011011011010011", 																																		
																	300 => "00000110001011110000011000101111", 301 => "00000011101100010000001110110001", 302 => "11100010111000001110001011100000", 303 => "00000100111010010000010011101001", 304 => "00000010010101100000001001010110", 305 =>"00000111110011000000011111001100", 306 => "01110111000000000111011100000000", 307 => "00000000101101000000000010110100", 308 => "00010110100000110001011010000011", 309 => "11111000100000111111100010000011", 310 => "01100000100001110110000010000111",311 => "01000101010000010100010101000001", 312 => "00100000000000000010000000000000", 313 => "01110101000001010111010100000101", 314 => "00010100000010110001010000001011", 315 => "01101000001010000110100000101000", 316 => "01010100000000100101010000000010"
																	,317 => "00000011001000000000001100100000", 318 => "00000000100011000000000010001100", 319 => "01000011010000000100001101000000", 320 => "00000110111010110000011011101011", 321 => "11000000011000001100000001100000", 322 => "00000001100001110000000110000111", 323 => "00001111001000000000111100100000", 324 => "00000000101110000000000010111000", 325 => "00000011000001000000001100000100", 326 => "01011001000001100101100100000110", 327 => "10100000110101011010000011010101"
																	,328 => "00000110101101110000011010110111", 329 =>"00000011010010110000001101001011", 330 => "11111101110000001111110111000000", 331 => "00000000100001000000000010000100", 332 => "00000001110000010000000111000001", 333 => "00000001000001110000000100000111", 334 => "11011000001000001101100000100000", 335 => "01010010010000010101001001000001", 336 => "11000001000101001100000100010100", 337 => "00100000100100010010000010010001", 338 => "01000100000100110100010000010011", 339 => "10100000101010111010000010101011"
																	,340 => "00000110000010010000011000001001", 341 => "00000001001101000000000100110100", 342 => "10000001001000001000000100100000", 343 => "00000111101011110000011110101111", 344 => "11000101000000001100010100000000", 345 => "00000011000111000000001100011100", 346 => "00000100101000000000010010100000", 347 => "10000100000010011000010000001001", 348 => "10000000000010101000000000001010", 349 => "10000011001010011000001100101001", 350 => "10000001000000001000000100000000", 351 => "00010010000011000001001000001100"
																	,352 => "00000000001100010000000000110001", 353 => "00000101000100010000010100010001", 354 => "10001110111000001000111011100000", 355 => "00000110111011010000011011101101", 356 =>"00000001111111110000000111111111", 357 => "00000000111001010000000011100101", 358 =>"11111001011000001111100101100000", 359 =>"11101110000011011110111000001101", 360 =>"00001010100000010000101010000001", 361 => "10000010010100101000001001010010", 362 => "01110000011110100111000001111010", 363 =>"00010011000001100001001100000110", 364 =>"01000100000110110100010000011011", 365 => "01101010000000000110101000000000"
																	,366 => "00000011100100010000001110010001", 367 => "00000101010011110000010101001111", 368 => "01111011101000000111101110100000", 369 => "00000010100011110000001010001111", 370 =>"00110101100000000011010110000000", 371 => "00000110010011010000011001001101", 372 =>"00011101010000000001110101000000", 373 => "11000000110000011100000011000001", 374 => "11101000001100001110100000110000", 375 => "00001000000010000000100000001000", 376 => "10110110000010001011011000001000", 377 =>"10010000010100111001000001010011", 378 =>"01110000010110100111000001011010"
																	,379 =>"00000100010001100000010001000110", 380 => "00000110011100100000011001110010", 381 =>"11000001000000001100000100000000", 382 =>"00000001111101010000000111110101", 383 =>"00000000001101000000000000110100", 384 => "00000010100110000000001010011000", 385 => "00100111111000000010011111100000", 386 => "11011001100000101101100110000010", 387 => "11000100000110001100010000011000", 388 => "01001001100000110100100110000011", 389 => "01000001001000010100000100100001", 390 => "01010000010100110101000001010011", 391 => "01101010110000010110101011000001", 392 => "10000100000110111000010000011011", 393 => "10100000000100101010000000010010", 394 => "10000010000000011000001000000001", 395 => "11100000110101011110000011010101", 396 => "00100100000110110010010000011011"
																	,397 => "01001101101010110100110110101011", 398 => "00000110011010010000011001101001", 399 => "00110010011000010011001001100001",																	
																	400 => "10111110001011111011111000101111", 401 => "10111011101100011011101110110001", 402 => "11100010111101111110001011110111", 403 => "10011101011110011001110101111001", 404 => "10101110101011001010111010101100", 405 =>"11111001011111001111100101111100", 406 => "01110111101110000111011110111000", 407 => "00010101111101000001010111110100", 408 => "00010110111101110001011011110111", 409 => "11011111110001111101111111000111", 410 => "01110001011101110111000101110111",411 => "01101110001010110110111000101011", 412 => "01011101000000000101110100000000", 413 => "01110101101111010111010110111101", 414 => "00010111010110110001011101011011", 415 => "01101011111010000110101111101000", 416 => "01010101011100100101010101110010"
																	,417 => "10111101100100001011110110010000", 418 => "01011100100011000101110010001100", 419 => "01001011100110100100101110011010", 420 => "11011101111010111101110111101011", 421 => "11011110000000111101111000000011", 422 => "00111011100001110011101110000111", 423 => "00101110011110010010111001111001", 424 => "00010111101110000001011110111000", 425 => "00001011100111000000101110011100", 426 => "01011010111011100101101011101110", 427 => "10111011110101011011101111010101"
																	,428 => "10111110101101111011111010110111", 429 =>"01101101110010110110110111001011", 430 => "11111101111011101111110111101110", 431 => "00010101110001000001010111000100", 432 => "10111011100100011011101110010001", 433 => "00100101110001110010010111000111", 434 => "11011010111000011101101011100001", 435 => "01010101110100110101010111010011", 436 => "11101011100101001110101110010100", 437 => "00110101110100010011010111010001", 438 => "01010111001100110101011100110011", 439 => "11011101101010111101110110101011"
																	,440 => "10111110000010011011111000001001", 441 => "00101011101101000010101110110100", 442 => "10010111000010011001011100001001", 443 => "11011111101011111101111110101111", 444 => "11000101011110001100010101111000", 445 => "01100101110111000110010111011100", 446 => "00010111001001010001011100100101", 447 => "10001011101100011000101110110001", 448 => "10001011100010101000101110001010", 449 => "11101011101010011110101110101001", 450 => "11000001011100001100000101110000", 451 => "01011100100111000101110010011100"
																	,452 => "10111000001100011011100000110001", 453 => "10100101110100011010010111010001", 454 => "10010111011101111001011101110111", 455 => "11011110111011011101111011101101", 456 =>"01111110111111110111111011111111", 457 => "10011100101111111001110010111111", 458 =>"11111010111010111111101011101011", 459 =>"11101111011111011110111101111101", 460 =>"00010111001010110001011100101011", 461 => "11001010101110101100101010111010", 462 => "01111111011110100111111101111010", 463 =>"00101110100111100010111010011110", 464 =>"01000111101110110100011110111011", 465 => "01011111010100000101111101010000"
																	,466 => "10111011100100011011101110010001", 467 => "10100101110100011010010111010001", 468 => "01110111110111010111011111011101", 469 => "01010101110011110101010111001111", 470 =>"00110110111011000011011011101100", 471 => "11001010111011011100101011101101", 472 =>"00101110111010100010111011101010", 473 => "11110101110000011111010111000001", 474 => "11101110111100001110111011110000", 475 => "00101110010010000010111001001000", 476 => "10101111101110001010111110111000", 477 =>"10101110110100111010111011010011", 478 =>"01111011101110100111101110111010"
																	,479 =>"10111100010001101011110001000110", 480 => "11001110111100101100111011110010", 481 =>"11000101110010001100010111001000", 482 =>"00111011111101010011101111110101", 483 =>"00001101011101000000110101110100", 484 => "01010101110110000101010111011000", 485 => "00100111101111110010011110111111", 486 => "11011010111011101101101011101110", 487 => "11010111001110001101011100111000", 488 => "01001011110011110100101111001111", 489 => "01110111001000010111011100100001", 490 => "01011110110100110101111011010011", 491 => "01110111010101110111011101010111", 492 => "10000101111110111000010111111011", 493 => "10100101110100101010010111010010", 494 => "10001011100100011000101110010001", 495 => "11111010111101011111101011110101", 496 => "00100101111110110010010111111011"
																	,497 => "10111110110101011011111011010101", 498 => "10111011001101001011101100110100", 499 => "10111001100100111011100110010011",																	
																	500 => "00111110001011110011111000101111", 501 => "01110100111100010111010011110001", 502 => "11100010011101111110001001110111", 503 => "10011001111010011001100111101001", 504 => "10010101001111001001010100111100", 505 =>"11100111110011001110011111001100", 506 => "00111011101110000011101110111000", 507 => "00111000101101000011100010110100", 508 => "00111000101101110011100010110111", 509 => "11001111110001111100111111000111", 510 => "01001111100001110100111110000111", 511 => "01000011101010110100001110101011", 512 => "00100011100000000010001110000000", 513 => "01110001111011010111000111101101", 514 => "00001110010110110000111001011011", 515 => "01001111011010000100111101101000", 516 => "01010100011100100101010001110010"
																	,517 => "00111011001000000011101100100000", 518 => "00010001110011000001000111001100", 519 => "01000111000110100100011100011010", 520 => "11011100111010111101110011101011", 521 => "11000000111000111100000011100011", 522 => "00001111100001110000111110000111", 523 => "00111000011110010011100001111001", 524 => "00111000101110000011100010111000", 525 => "00111000000111000011100000011100", 526 => "00011110110011100001111011001110", 527 => "10011101110101011001110111010101"
																	,528 => "00111110101101110011111010110111", 529 =>"01100011110010110110001111001011", 530 => "11111001111011101111100111101110", 531 => "00010011100001000001001110000100", 532 => "01110010000111010111001000011101", 533 => "00011101000001110001110100000111", 534 => "00111110110000010011111011000001", 535 => "00011110100100110001111010010011", 536 => "00111111000101000011111100010100", 537 => "00011101100100010001110110010001", 538 => "01001110001100110100111000110011", 539 => "10100111101010111010011110101011"
																	,540 => "00111110000010010011111000001001", 541 => "00100110011101000010011001110100", 542 => "10000001110010011000000111001001", 543 => "11110001111011111111000111101111", 544 => "11000101000011101100010100001110", 545 => "00011111000111000001111100011100", 546 => "00111000001001010011100000100101", 547 => "00111100001100010011110000110001", 548 => "00111100000010100011110000001010", 549 => "00111111001010010011111100101001", 550 => "11001110000000001100111000000000", 551 => "00000111100111000000011110011100"
																	,552 => "00111000001100010011100000110001", 553 => "10100000111100011010000011110001", 554 => "10000011111101111000001111110111", 555 => "11000111111011011100011111101101", 556 =>"01111110011111110111111001111111", 557 => "10011100111001011001110011100101", 558 =>"00111111110010110011111111001011", 559 =>"11001111011111011100111101111101", 560 =>"00111000001010110011100000101011", 561 => "11001110010100101100111001010010", 562 => "00111011111110100011101111111010", 563 =>"00000111100111100000011110011110", 564 =>"01000011101110110100001110111011", 565 => "01100011110100000110001111010000"
																	,566 => "00111011100100010011101110010001", 567 => "10101001100111111010100110011111", 568 => "01110011110111010111001111011101", 569 => "01010001110011110101000111001111", 570 =>"00110100011111000011010001111100", 571 => "11001110010011011100111001001101", 572 =>"00111000111010100011100011101010", 573 => "00111111100000010011111110000001", 574 => "00111111011100000011111101110000", 575 => "00111000010010000011100001001000", 576 => "10011101101110001001110110111000", 577 =>"10011010001110111001101000111011", 578 =>"01001111110110100100111111011010"
																	,579 =>"00111100010001100011110001000110", 580 => "11001100111100101100110011110010", 581 =>"11000000111010001100000011101000", 582 =>"00111110001111010011111000111101", 583 =>"00001100100001110000110010000111", 584 => "01010011100110000101001110011000", 585 => "00111001001111110011100100111111", 586 => "10011110110011101001111011001110", 587 => "00111110001110000011111000111000", 588 => "00111010010011110011101001001111", 589 => "00111011001000010011101100100001", 590 => "00011110110100110001111011010011", 591 => "01100111010101110110011101010111", 592 => "10000001111110111000000111111011", 593 => "10100001110100101010000111010010", 594 => "10000111000100011000011100010001", 595 => "11111000111101011111100011110101", 596 => "00100111001110110010011100111011"
																	,597 => "00111110110101010011111011010101", 598 => "01100100111101000110010011110100", 599 => "00110010011111110011001001111111",																	
														      	600 => "01011110001011110101111000101111", 601 => "01011011101100010101101110110001", 602 => "01011111000101110101111100010111", 603 => "01011100111010010101110011101001", 604 => "01011100101011000101110010101100", 605 =>"01011111110011000101111111001100", 606 => "01011011101110000101101110111000", 607 => "01011000101101000101100010110100", 608 => "01011000101101110101100010110111", 609 => "01011111110001110101111111000111", 610 => "01011011100001110101101110000111",611 => "01011010001010110101101000101011", 612 => "01011001000000000101100100000000", 613 => "01011011101011010101101110101101", 614 => "01011000010110110101100001011011", 615 => "01011011011010000101101101101000", 616 => "01011010101000100101101010100010"
																	,617 => "01011011001000000101101100100000", 618 => "01011000100011000101100010001100", 619 => "01011010000110100101101000011010", 620 => "01011110111010110101111011101011", 621 => "01011110000000110101111000000011", 622 => "01011001100001110101100110000111", 623 => "01011000011110010101100001111001", 624 => "01011000101110000101100010111000", 625 => "01011000000111000101100000011100", 626 => "01011010110011100101101011001110", 627 => "01011101110101010101110111010101"
																	,628 => "01011110101101110101111010110111", 629 =>"01011011010010110101101101001011", 630 => "01011111111011100101111111101110", 631 => "01011000100001000101100010000100", 632 => "01011011100100010101101110010001", 633 => "01011001000001110101100100000111", 634 => "01011110110000010101111011000001", 635 => "01001011100100110100101110010011", 636 => "01011111000101000101111100010100", 637 => "01011001100100010101100110010001", 638 => "01011010001100110101101000110011", 639 => "01011101101010110101110110101011"
																	,640 => "01011110000010010101111000001001", 641 => "01011001001101000101100100110100", 642 => "01011100000010010101110000001001", 643 => "01011111101011110101111110101111", 644 => "01011110001010000101111000101000", 645 => "01011011000111000101101100011100", 646 => "01011000001001010101100000100101", 647 => "10010110001100011001011000110001", 648 => "01011100000010100101110000001010", 649 => "01011111001010010101111100101001", 650 => "01011110000000000101111000000000", 651 => "01011000100111000101100010011100"
																	,652 => "00000110001111110000011000111111", 653 => "01011101000100010101110100010001", 654 => "01011100011101110101110001110111", 655 => "01011110111011010101111011101101", 656 =>"01011011111111110101101111111111", 657 => "01011100111001010101110011100101", 658 =>"01011111110010110101111111001011", 659 =>"01011111011111010101111101111101", 660 =>"01011000001010110101100000101011", 661 => "01011110010100100101111001010010", 662 => "01011011111110100101101111111010", 663 =>"01011000100111100101100010011110", 664 =>"01011010001110110101101000111011", 665 => "01011011010100000101101101010000"
																	,666 => "01011011100100010101101110010001", 667 => "01011101010011110101110101001111", 668 => "01011011110111010101101111011101", 669 => "01011010100011110101101010001111", 670 =>"01011001101011000101100110101100", 671 => "01011110010011010101111001001101", 672 =>"01011000111010100101100011101010", 673 => "01011111100000010101111110000001", 674 => "01011111011100000101111101110000", 675 => "01011000010010000101100001001000", 676 => "01011101101110000101110110111000", 677 =>"01011100110100110101110011010011", 678 =>"01011011110110100101101111011010"
																	,679 =>"01011100010001100101110001000110", 680 => "01011110011100100101111001110010", 681 =>"10101110000010001010111000001000", 682 =>"01011001111101010101100111110101", 683 =>"01011000011001000101100001100100", 684 => "01011010100110000101101010011000", 685 => "01011001001111110101100100111111", 686 => "01011110110011100101111011001110", 687 => "01011110001110000101111000111000", 688 => "01011010010011110101101001001111", 689 => "01011011001000010101101100100001", 690 => "01011010110100110101101011010011", 691 => "01011011010101110101101101010111", 692 => "01011100001110110101110000111011", 693 => "01011101000100100101110100010010", 694 => "01011100000100010101110000010001", 695 => "01011111110101010101111111010101", 696 => "01011001001110110101100100111011"
																	,697 => "01011110110101010101111011010101", 698 => "01011011001101000101101100110100", 699 => "01011001100100110101100110010011",																	
												    				700 => "10010110001011111001011000101111", 701 => "10010011101100011001001110110001", 702 => "10010111000101111001011100010111", 703 => "10010100111010011001010011101001", 704 => "10010100101011001001010010101100", 705 =>"10010111110011001001011111001100", 706 => "10010011101110001001001110111000", 707 => "10010000101101001001000010110100", 708 => "10010000101101111001000010110111", 709 => "10010111110001111001011111000111", 710 => "10010011100001111001001110000111",711 => "10010010001010111001001000101011", 712 => "10010001000000001001000100000000", 713 => "10010011101011011001001110101101", 714 => "10010000010110111001000001011011", 715 => "10010011011010001001001101101000", 716 => "10010010101000101001001010100010"
																	,717 => "10010011001000001001001100100000", 718 => "10010000100011001001000010001100", 719 => "10010010000110101001001000011010", 720 => "10010110111010111001011011101011", 721 => "10010110000000111001011000000011", 722 => "10010001100001111001000110000111", 723 => "10010000011110011001000001111001", 724 => "10010000101110001001000010111000", 725 => "10010000000111001001000000011100", 726 => "10010010110011101001001011001110", 727 => "10010101110101011001010111010101"
																	,728 => "10010110101101111001011010110111", 729 =>"10010011010010111001001101001011", 730 => "10010111111011101001011111101110", 731 => "10010000100001001001000010000100", 732 => "10010011100100011001001110010001", 733 => "10010001000001111001000100000111", 734 => "10010110110000011001011011000001", 735 => "10010010100100111001001010010011", 736 => "10010111000101001001011100010100", 737 => "10010001100100011001000110010001", 738 => "10010010001100111001001000110011", 739 => "10010101101010111001010110101011"
																	,740 => "10010110000010011001011000001001", 741 => "10010001001101001001000100110100", 742 => "10010100000010011001010000001001", 743 => "10010111101011111001011110101111", 744 => "10010110001010001001011000101000", 745 => "10010011000111001001001100011100", 746 => "10010000001001011001000000100101", 747 => "10010100001100011001010000110001", 748 => "10010100000010101001010000001010", 749 => "10010111001010011001011100101001", 750 => "10010110000000001001011000000000", 751 => "10010000100111001001000010011100"
																	,752 => "10010000001100011001000000110001", 753 => "10010101000100011001010100010001", 754 => "10010100011101111001010001110111", 755 => "10010110111011011001011011101101", 756 =>"10010011111111111001001111111111", 757 => "10010100111001011001010011100101", 758 =>"10010111110010111001011111001011", 759 =>"10010111011111011001011101111101", 760 =>"10010000001010111001000000101011", 761 => "10010110010100101001011001010010", 762 => "10010011111110101001001111111010", 763 =>"10010000100111101001000010011110", 764 =>"10010010001110111001001000111011", 765 => "10010011010100001001001101010000"
																	,766 => "10010011100100011001001110010001", 767 => "10010101010011111001010101001111", 768 => "10010011110111011001001111011101", 769 => "10010010100011111001001010001111", 770 =>"10010001101011001001000110101100", 771 => "10010110010011011001011001001101", 772 =>"10010000111010101001000011101010", 773 => "10010111100000011001011110000001", 774 => "10010111011100001001011101110000", 775 => "10010000010010001001000001001000", 776 => "10010101101110001001010110111000", 777 =>"10010100110100111001010011010011", 778 =>"10010011110110101001001111011010"
																	,779 =>"10010100010001101001010001000110", 780 => "10010110011100101001011001110010", 781 =>"10010110000010001001011000001000", 782 =>"10010001111101011001000111110101", 783 =>"10010000011001001001000001100100", 784 => "10010010100110001001001010011000", 785 => "10010001001111111001000100111111", 786 => "10010110110011101001011011001110", 787 => "10010110001110001001011000111000", 788 => "10010010010011111001001001001111", 789 => "10010011001000011001001100100001", 790 => "10010010110100111001001011010011", 791 => "10010011010101111001001101010111", 792 => "10010100001110111001010000111011", 793 => "10010101000100101001010100010010", 794 => "10010100000100011001010000010001", 795 => "10010111110101011001011111010101", 796 => "10010001001110111001000100111011"
																	,797 => "10010110110101011001011011010101", 798 => "10010011001101001001001100110100", 799 => "10010001100100111001000110010011",																
																	800 => "10010110001011111001011000101111", 801 => "10010011101100011001001110110001", 802 => "11001011000101111100101100010111", 803 => "10010100111010011001010011101001", 804 => "10010100101011001001010010101100", 805 =>"10010111110011001001011111001100", 806 => "10010011101110001001001110111000", 807 => "10010000101101001001000010110100", 808 => "10010000101101111001000010110111", 809 => "10010111110001111001011111000111", 810 => "10010011100001111001001110000111",811 => "10010010001010111001001000101011", 812 => "10010001000000001001000100000000", 813 => "10010011101011011001001110101101", 814 => "10010000010110111001000001011011", 815 => "10010011011010001001001101101000", 816 => "10010010101000101001001010100010"
																	,817 => "10010011001000001001001100100000", 818 => "10010000100011001001000010001100", 819 => "10010010000110101001001000011010", 820 => "10010110111010111001011011101011", 821 => "10010110000000111001011000000011", 822 => "10010001100001111001000110000111", 823 => "10010000011110011001000001111001", 824 => "10010000101110001001000010111000", 825 => "10010000000111001001000000011100", 826 => "10010010110011101001001011001110", 827 => "10010101110101011001010111010101"
																	,828 => "10010110101101111001011010110111", 829 =>"10010011010010111001001101001011", 830 => "10010111111011101001011111101110", 831 => "10010000100001001001000010000100", 832 => "10010011100100011001001110010001", 833 => "10010001000001111001000100000111", 834 => "10010110110000011001011011000001", 835 => "10010010100100111001001010010011", 836 => "10010111000101001001011100010100", 837 => "10010001100100011001000110010001", 838 => "10010010001100111001001000110011", 839 => "10010101101010111001010110101011"
																	,840 => "10010110000010011001011000001001", 841 => "10010001001101001001000100110100", 842 => "10010100000010011001010000001001", 843 => "10010111101011111001011110101111", 844 => "10010110001010001001011000101000", 845 => "10010011000111001001001100011100", 846 => "10010000001001011001000000100101", 847 => "10010100001100011001010000110001", 848 => "10010100000010101001010000001010", 849 => "10010111001010011001011100101001", 850 => "10010110000000001001011000000000", 851 => "10010000100111001001000010011100"
																	,852 => "10010000001100011001000000110001", 853 => "10010101000100011001010100010001", 854 => "10010100011101111001010001110111", 855 => "10010110111011011001011011101101", 856 =>"10010011111111111001001111111111", 857 => "10010100111001011001010011100101", 858 =>"10010111110010111001011111001011", 859 =>"10010111011111011001011101111101", 860 =>"10010000001010111001000000101011", 861 => "10010110010100101001011001010010", 862 => "10010011111110101001001111111010", 863 =>"10010000100111101001000010011110", 864 =>"10010010001110111001001000111011", 865 => "10010011010100001001001101010000"
																	,866 => "10010011100100011001001110010001", 867 => "10010101010011111001010101001111", 868 => "10010011110111011001001111011101", 869 => "10010010100011111001001010001111", 870 =>"10010001101011001001000110101100", 871 => "10010110010011011001011001001101", 872 =>"10010000111010101001000011101010", 873 => "10010111100000011001011110000001", 874 => "10010111011100001001011101110000", 875 => "10010000010010001001000001001000", 876 => "10010101101110001001010110111000", 877 =>"10010100110100111001010011010011", 878 =>"10010011110110101001001111011010"
																	,879 =>"10010100010001101001010001000110", 880 => "10010110011100101001011001110010", 881 =>"10010110000010001001011000001000", 882 =>"10010001111101011001000111110101", 883 =>"10010000011001001001000001100100", 884 => "10010010100110001001001010011000", 885 => "10010001001111111001000100111111", 886 => "10010110110011101001011011001110", 887 => "10010110001110001001011000111000", 888 => "10010010010011111001001001001111", 889 => "10010011001000011001001100100001", 890 => "10010010110100111001001011010011", 891 => "10010011010101111001001101010111", 892 => "10010100001110111001010000111011", 893 => "10010101000100101001010100010010", 894 => "10010100000100011001010000010001", 895 => "10010111110101011001011111010101", 896 => "10010001001110111001000100111011"
																	,897 => "10010110110101011001011011010101", 898 => "10010011001101001001001100110100", 899 => "10010001100100111001000110010011",
																	900 => "00001110001011110000111000101111", 901 => "01110110001000010111011000100001", 902 => "11100010111000011110001011100001", 903 => "10011101001000011001110100100001", 904 => "10010101100000011001010110000001", 905 =>"00001111110011000000111111001100", 906 => "01110111000000010111011100000001", 907 => "00010110100000010001011010000001", 908 => "00001000101101110000100010110111", 909 => "11100001110001111110000111000111", 910 => "00001011100001110000101110000111",911 => "00001010001010110000101000101011", 912 => "00000101000000000000010100000000", 913 => "00001011101011010000101110101101", 914 => "00001000010110110000100001011011", 915 => "00001011011010000000101101101000", 916 => "00001010101000100000101010100010"
																	,917 => "00001011001000000000101100100000", 918 => "00010001100000010001000110000001", 919 => "11100010111000011110001011100001", 920 => "11011101011000011101110101100001", 921 => "11000000011000011100000001100001", 922 => "00001001100001110000100110000111", 923 => "00001111001000010000111100100001", 924 => "00010111000000010001011100000001", 925 => "00001000000111000000100000011100", 926 => "01000010110011100100001011001110", 927 => "10000101110101011000010111010101"
																	,928 => "00001110101101110000111010110111", 929 =>"01101001011000010110100101100001", 930 => "11111101110000011111110111000001", 931 => "00010000100000010001000010000001", 932 => "01110010001000010111001000100001", 933 => "00001001000001110000100100000111", 934 => "11011000001000011101100000100001", 935 => "01010010011000010101001001100001", 936 => "00001111000101000000111100010100", 937 => "00000101100100010000010110010001", 938 => "00001010001100110000101000110011", 939 => "00001101101010110000110110101011"
																	,940 => "00001110000010010000111000001001", 941 => "00100110100000010010011010000001", 942 => "10000001001000011000000100100001", 943 => "11110101111000011111010111100001", 944 => "11000101000000011100010100000001", 945 => "00001011000111000000101100011100", 946 => "00000100101000010000010010100001", 947 => "10000110001000011000011000100001", 948 => "00001100000010100000110000001010", 949 => "00001111001010010000111100101001", 950 => "00001110000000000000111000000000", 951 => "00001000100111000000100010011100"
																	,952 => "00001000001100010000100000110001", 953 => "10100010001000011010001000100001", 954 => "10001110111000011000111011100001", 955 => "11011101101000011101110110100001", 956 =>"01111111111000010111111111100001", 957 => "00001100111001010000110011100101", 958 =>"11111001011000011111100101100001", 959 =>"11101111101000011110111110100001", 960 =>"00001000001010110000100000101011", 961 => "00001110010100100000111001010010", 962 => "00001011111110100000101111111010", 963 =>"00001000100111100000100010011110", 964 =>"01000010001110110100001000111011", 965 => "00001011010100000000101101010000"
																	,966 => "00001011100100010000101110010001", 967 => "10101001111000011010100111100001", 968 => "01111011101000010111101110100001", 969 => "01010001111000010101000111100001", 970 =>"00110101100000010011010110000001", 971 => "00001110010011010000111001001101", 972 =>"00011101010000010001110101000001", 973 => "11110000001000011111000000100001", 974 => "00001111011100000000111101110000", 975 => "00001000010010000000100001001000", 976 => "00001101101110000000110110111000", 977 =>"00001100110100110000110011010011", 978 =>"00000111110110100000011111011010"
																	,979 =>"00001100010001100000110001000110", 980 => "11001110010000011100111001000001", 981 =>"11000001000000011100000100000001", 982 =>"00111110101000010011111010100001", 983 =>"00001100100000010000110010000001", 984 => "00001010100110000000101010011000", 985 => "00100111111000010010011111100001", 986 => "11011001110000011101100111000001", 987 => "00001110001110000000111000111000", 988 => "00001010010011110000101001001111", 989 => "00001011001000010000101100100001", 990 => "00001010110100110000101011010011", 991 => "00000111010101110000011101010111", 992 => "00001100001110110000110000111011", 993 => "00001101000100100000110100010010", 994 => "00001100000100010000110000010001", 995 => "00001111110101010000111111010101", 996 => "00001001001110110000100100111011"
																	,997 => "00001110110101010000111011010101", 998 => "01100110100000010110011010000001", 999 => "00110010011000010011001001100001"
																	);
																	
																	
																																												-------------------------------
																	
	signal DataOutput2 : DataTypeOutput := (0 => "11111110110111110111111011011111", 1 => "11111100101111011111110010111100", 2 => "11111101011001101111110101101100",3 => "11111111101110101111111110111000", 4 => "11111111100110111101111110011011"
																	,5 => "11111001100111111101100110011011",6 => "10000010111111101000001011101110", 7 => "01100111111011100110110111101110", 8 => "11101111111110111110101111111011", 9 => "10010111001111101001011100111111",10 => "11111100111111111111110011111110",
																	11 => "11111001100111111101100110010111", 12 => "11110001111111011111000110111101",13 => "11110011111001111101101111100111",14 => "11110000010001001110000001000100",15 => "11110010101011111111001010101100",16 => "11110010000111010111001000011100",
																	17 => "11111000000011111101100000000111",18 => "11110000111010001111000011001000",19 => "11110000000111101110010000011110", 20 => "11110001011011111110000101101111",21 => "11110010010011011111001001001110",22 => "11110010010110100111001001011010", 23 => "11110011100100111101001110010011"
																	,24 => "11110011000110011011001100001001", 25 => "00000110000111110000011010011111", 26 => "00000110100110101010011010011010", 27 => "00000000001110101000000000111010", 28 => "00000100110111000000010011101100", 29 => "00000000111101010000000011100101", 30 => "00000001111110010000000111111101", 31 => "00000111001000010000011100000001"
																   ,32 => "11111011110100111011101111000011",33 => "10110111111001111011011110100111",34 => "10110011111010001001101111101000",35 => "10101101101111111011110110111111",36 => "10111111101101001011111110110111",37 => "01111101111101111111110111110111",38 => "10111110001101101001111001101101"
																	,39 => "11111010011111111011101001101111",40 => "10011111100011011001111111001101",41 => "10111110011101111001011001110111" ,42 => "00110111111000100001011111100010",43 => "00100101111111010010010111111011",44 =>"10110011111010100011001111101010", 45 =>"10101110111111011000111011111101",46 =>"11101001111100101100100111110010"
																	,47 => "11111100001110011011110000101001", 48 => "10101111110010001010111101001000", 49 => "01111101111110101101110111111010", 50 => "01011111101110001101111110111000", 51 => "11011101110111111101110111101111", 52 =>"01101101111100100110110111111010",53 => "00111111111111100011111111111100"
																	,54 => "11111100100011011011110010001101",55 => "11111111111110111111111110111011",56 => "10111111010100101001011101010010",57 => "00011111110100100000111111010010", 58 => "00011111111001100001111111100000", 59 => "11111110100010001111111010001010", 60 => "11111101111100011111110111110000"
																	,61 => "11111011000011111011101100001111", 62 => "00111001111101010011100101110101", 63 => "11011011100111110111101110011111", 64 => "11110101111111101111010111111110", 65 => "11110111110110101111011111101010", 66 => "11111110101111111111111010101111", 67 => "01101111111011110110111111100111"
																	,68 => "11111000100111001011100010011100",69 => "11110011111110101011001110111010", 70 => "00111111001111100110111100111110", 71 => "11001011001110111000101100111011", 72 => "00111110011001000011111001111100", 73 => "10011110011101011001111001111101", 74 => "11100000110010001110000011001100"
																	,75 => "00110011010010110011001101101011",76 => "00001111011110100100111101111010", 77 => "00011100111000000100110011100000", 78 => "10000000111001101100000011100110", 79 => "01011111001010000101111100110000", 80 => "11001111001100111100111100111011", 81 => "11011000000100101101100000010110"
																	,82 => "11010000100010001101000010011000",83 => "00101101101011000110110110101100", 84 => "10000111001110011101011100111001", 85 => "00100110011000010110011001100001", 86 => "01011010011110100101101001100010", 87 => "01111011110001110111101111001111", 88 => "01101111001111010110111100111001"
																	,89 => "11010111001011001101011100111100", 90 => "00100111001110001010011100111000", 91 => "11110011100110110101001110011011", 92 => "11101001110111000110100111011100", 93 => "01011100110000010101110011110001", 94 => "01111001100001000111100110010100", 95 =>"00110011000011000011001100001000"
																	,96 => "01101101100011100110110110011110", 97 => "01001001100000011100100110000001", 98 => "00001001100001111010100110000111",99 => "01111100111000010011110011100001",																	
																	100 => "10000001100011101000000110011110", 101 => "10111100111101111011110011110110", 102 => "00110011000100011011001100010011"
																	,103 => "10101101110011011010110111001111",104 => "10010011100111101001001110011100",105 => "00101111100111000110111110011101",106 => "10011100110101001001110011010101", 107 => "11101010011010101110111001111010", 108 => "01111011100111110101101110011111", 109 => "00011010100110100101101010011010",
																	110 => "01000100010101000100011001010100",111 => "11010101010101001101010101010101", 112 => "00010011101010110101001110101010",113 => "11010101101110011101010110111000", 114 => "11010001100110001101010110001000", 115 => "10010011101010011011001110101001", 116 =>"10110101010100101001010101010010",
																	117 => "01010000110111110101001011011111", 118 => "10111000011110011011100001111111", 119 => "01010001100111011101000110011111", 120 => "11101010100101011110101010010001", 121 => "10111010100110101010101011011010", 122 => "10101001101011010010100110101101", 123 => "11101010111101101110101011110111", 124 => "11010101010101011111010101010101", 125 => "00101101010101000010110100010100", 126 => "01011101010111101101110101011110", 127 => "10010100110100101001110011010010", 128 => "00101010011000101010101001100010", 129 => "10001011001001001010101100100100", 130 => "11000010101101011100001010100101", 131 => "10010101000111111001010100011101"
																	,132 => "10010001000010101001010100001010", 133 => "01101001001011000110100100101000", 134 => "01110101111100100111010111110111", 135 => "10100110100111011010011010010101", 136 => "10000111011011001010011111101100", 137 => "00101100000101010010110000010100", 138 => "01010100101010100101010010101000", 139 => "00101100001010100110110000101010", 140 => "00011110110101010001111001010101", 141 => "11011011010101011101101101010100", 142 =>"11011010101001011101001010100101", 143 => "01101101010101001110110101010100"
																	,144 => "00001000100010000000101010001000", 145 => "11011101010111111101110101010111", 146 => "11010101001100011101010100110100", 147 => "10101010110000111010101011001011", 148 => "10001011011000001010101111100000", 149 => "00101010010010010010101001001000", 150 =>"10101101010111111010110101011110", 151 => "10010011010101111011001101010111", 152 =>"00110110010101000011011001110100", 153 => "10001101010101101100110101010110", 154 => "01001010100110110100111010011011", 155 => "10110110101010111111011010101011", 156 => "10101010100010101011101010001010", 157 => "10101001010111101010100101010110", 158 => "00101010011100110010101001110010", 159 => "11101010111001111110101011100011"
																	,160 => "01010001100111110101001110011111",161 => "10111010101010101011101010101000", 162 => "00110101010100111011010101010001", 163 => "11010101101101101101010110110010", 164 => "10111010010000101010101000000010", 165 => "00100101010001001010010101000100", 166 => "01110101010101010111010101010100", 167 => "01111010101110000101101010111000", 168 => "00101000101010010010100011101001", 169 => "10010101101010100001010110101010", 170 => "01100110101010100110111010101010", 171 => "11011100101010010101110010101001", 172 => "10101001100011101000100110001110", 173 => "10101001011110111010100101101011", 174 => "11101010111001001110101011100110", 175 => "11101010110110011110101011010001", 176 => "10001010101000111000101010000011", 177 => "01010100110101100101010011110110", 178 => "01011101010111010101010101011101", 179 => "11101101110101100110110111010111", 180 => "00101001010110011010100101011000", 181 => "01110101011111100111010101100110"
																	,182 => "01010001101010110101010110101011", 183 => "00101001010101000010100101010000", 184 => "11011010101011101101101010101011", 185 => "10101110101000011010111010101001", 186 => "10001001101000111010100100100011", 187 => "01000110101011110100011010101110", 188 => "10110101010101001011010101010110", 189 => "01010101010100110001010101010011", 190 => "00101110101011100010111000101110", 191 => "11100100110101001110010011010101", 192 => "10101011001010101011101100101010", 193 => "00100110101001100010011010100111"
																	,194 => "11011010010111111101111001011111", 195 => "10110101010011011011010101001001", 196 => "10101010010111011010101001011000", 197 => "00001110101001110000111010101111", 198 => "10001010111010111010101001101011", 199 => "11010101010010011101010101001000", 																	
																	200 => "11000100101010111100010110101011", 201 => "01110101010111110111010101011001", 202 => "11101010100101010110101010010111", 203 => "10011010101011011001101010101001", 204 => "10000101111010101001010110101010", 205 =>"11101010110011001010101011001100", 206 => "10101001110110000010100111011000", 207 => "10101000101101001011101010110100", 208 =>"00101010010101100010101001010111", 209 => "11110101010001101111010101000111", 210 => "01110101010000110111011101000011", 211 => "01010101001010110111010100101011", 212 => "00100001010100000010100101010000", 213 => "01110101101011100111010110101010", 214 => "00010110101010111001011010101011", 215 => "01101010101101010110101010110100", 216 => "01010100101110100101010010101010"
																	,217 => "01100000101010000110010010101000", 218 => "00100110110111000010011011001100", 219 => "01011011000111110101101100011010", 220 => "11011101101101111101110110110101", 221 => "11100011111000111100001101100011", 222 => "00110011011001100011001101100111", 223 => "00011110110110110001111011011001", 224 => "00010111011010000101111101101000", 225 => "00011011000101000001101100011100", 226 => "01011011011011100101101101100110", 227 => "10111011010101011010101101010101"
																	,228 => "11010010111011111101011011101111", 229 =>"01101001011111100110100101110110", 230 => "11111011011011000111101101101110", 231 => "11011000100001011101100010000100", 232 => "01100110110100010111011010010001", 233 => "11011000100001110101100010000111", 234 => "11011011011000001101101101100001", 235 => "11011001010100111111110101010011", 236 => "11100101001100101110010100110110", 237 => "11011001100101011101100110010001", 238 => "01000110011101100100111001110110", 239 => "10110101011101111011010101110110"
																	,240 => "11000000001110111100000100111011", 241 => "11011001001111001101100100110100", 242 => "10101100000011001010110000001001", 243 => "11110101111011111111010111101101", 244 => "11111011101010001101101100101000", 245 => "01100011110110010110001111011000", 246 => "00001001011101000000100101110110", 247 => "10000110011101101100111001110110", 248 => "11011010000000101101101000001010", 249 => "11101010011111101110101001110110", 250 => "11011011000000001100101100000000", 251 => "11011000100111101101100010011100"
																	,252 => "00000100001110110000011000111011", 253 => "11011010100110011101101010001001", 254 => "10011101111010001001110111101101", 255 => "11011101101101111101110110110101", 256 =>"11001001101111111101100111111111", 257 => "11011010011001010101101001100101", 258 =>"11011011110010110101101111001011", 259 =>"11011011101111011101001010111101", 260 =>"11011000001010110101100000101011", 261 => "11011011010100100101101101010010", 262 => "11011001111110101101100011111010", 263 =>"11011000010011101100100001001110", 264 =>"11011001001110111101110100111011", 265 => "11011001101010011101100110101000"
																	,266 => "01110000001011110111001000101111", 267 => "11011010101101111101101010100111", 268 => "01111011010110000111101101011101", 269 => "01010011011001010101001101100111", 270 =>"11001001111011001101100110101100", 271 => "11011011010011010101101101001101", 272 =>"11011000111010100101100011101010", 273 => "11011011110000011100100111000001", 274 => "11011011011100101101101101110000", 275 => "11011000010010101101100001001000", 276 => "11011010110110001101111011011000", 277 =>"11011010011010111001101001101011", 278 =>"11011001110110101100100111011010"
																	,279 =>"10001000010110111000100011011011", 280 => "11110110001110101111011000110010", 281 =>"11000010110110011000001011011000", 282 =>"00111011011101010111101101110101", 283 =>"11011010011011001101100001100100", 284 => "11011001010110001100100101011000", 285 => "11011000100111111111100010011111", 286 => "11011011011001101101111111100110", 287 => "11011010001110000101101000111000", 288 => "11011000010011110101100001001111", 289 => "11011001100100011101100010010001", 290 => "11011001011010111111100101101011", 291 => "11011001101010111100100110101011", 292 => "10000111011100101000011101110110", 293 => "10100100101101101110010010110110", 294 => "10000100011101101010010001110110", 295 => "11110101011111101111010101110110", 296 => "00100111011101100010011101010110"
																	,297 => "11011000101110111101101010111011", 298 => "01100110111110100110011011011010", 299 => "00110110110101100011011011010011", 																																		
																	300 => "00000100001011110000011000101111", 301 => "00000011111100010000001110110001", 302 => "11100010111000100110001011100000", 303 => "00000100111010000000010011101001", 304 => "00010010000101100000001001010110", 305 =>"00000111110011000000010111001100", 306 => "01110111000001010111011100000000", 307 => "00000000101101000000001010110100", 308 => "00010110100000110011011010000011", 309 => "11111000100000101111100010000011", 310 => "01100000100001110110001010000111",311 => "01000101010000011100010101000001", 312 => "00100000001000000010000000000000", 313 => "01110101000011010111010100000101", 314 => "00010100000010111001010000001011", 315 => "01101000001010100110100000101000", 316 => "01010100000100100101010000000010"
																	,317 => "00000010001000000000001100100000", 318 => "00000000110011000000000010001100", 319 => "01000011010001010100001101000000", 320 => "00000110111010010000011011101011", 321 => "11100000111000001100000001100000", 322 => "00000001100001110000100110000111", 323 => "00001111001101000000111100100000", 324 => "00000000101110000000100010111000", 325 => "00000011000001001000001100000100", 326 => "01011001000000100101100100000110", 327 => "10100000110101011010100011010101"
																	,328 => "00000100101101110000011010110111", 329 =>"00000011011010110000001101001011", 330 => "11111101110000100111110111000000", 331 => "00000000100001010000000010000100", 332 => "00010001100000010000000111000001", 333 => "00000001000001110000010100000111", 334 => "11011000001010101101100000100000", 335 => "01010010010000010101011001000001", 336 => "11000001000101001000000100010100", 337 => "00100000100100110010000010010001", 338 => "01000100000100110100000000010011", 339 => "10100000101010101010000010101011"
																	,340 => "00000100000010010000011000001001", 341 => "00000001011101000000000100110100", 342 => "10000001001001011000000100100000", 343 => "00000111101011010000011110101111", 344 => "11100101100000001100010100000000", 345 => "00000011000111000000101100011100", 346 => "00000100101101000000010010100000", 347 => "10000100000010011000110000001001", 348 => "10000000000010100000000000001010", 349 => "10000011001011011000001100101001", 350 => "10000001000000001000100100000000", 351 => "00010010000011100001001000001100"
																	,352 => "00000000000100010000000000110001", 353 => "00000101001100010000010100010001", 354 => "10001110111001011000111011100000", 355 => "00000110111011110000011011101101", 356 =>"00010001101111110000000111111111", 357 => "00000000111001010000010011100101", 358 =>"11111001011001011111100101100000", 359 =>"11101110000011011110111100001101", 360 =>"00001010100000010000001010000001", 361 => "10000010010100101100001001010010", 362 => "01110000011110100111000011111010", 363 =>"00010011000001100000001100000110", 364 =>"01000100000110110100010010011011", 365 => "01101010000100000110101000000000"
																	,366 => "00000011100000010000001110010001", 367 => "00000101010111110000010101001111", 368 => "01111011101001010111101110100000", 369 => "00000010100011010000001010001111", 370 =>"00100101110000000011010110000000", 371 => "00000110010011010000001001001101", 372 =>"00011101010001010001110101000000", 373 => "11000000110000011100001011000001", 374 => "11101000001100001100100000110000", 375 => "00001000000010010000100000001000", 376 => "10110110000010001011010000001000", 377 =>"10010000010100111101000001010011", 378 =>"01110000010110100111001001011010"
																	,379 =>"00000100010000100000010001000110", 380 => "00000110011110100000011001110010", 381 =>"11000001000000011000000100000000", 382 =>"00000001111101010100000111110101", 383 =>"00000010001111000000000000110100", 384 => "00000010100110000000001000011000", 385 => "00100111111000010110011111100000", 386 => "11011001100000101101100100000010", 387 => "11000100000110001100110000011000", 388 => "01001001100000110000100110000011", 389 => "01000001001000010100000110100001", 390 => "01010000010100110111000001010011", 391 => "01101010110000010110101111000001", 392 => "10000100100110111000010000011011", 393 => "10100000000100101110000000010010", 394 => "10000010000100011000001000000001", 395 => "11100000110111011110000011010101", 396 => "00100100000110110010010010011011"
																	,397 => "01001101101000110100110110101011", 398 => "00000110011110010000011001101001", 399 => "00110010011001000011001001100001",																	
																	400 => "10111110001010111011111000101111", 401 => "10111011101110011011101110110001", 402 => "11100010111101010110001011110111", 403 => "10011101011110001001110101111001", 404 => "10111110111011001010111010101100", 405 =>"11111001011111101111100100111100", 406 => "01110111101110000111011110111000", 407 => "00010101111101000001010110110100", 408 => "00010110111101110101011011110111", 409 => "11011111110001011101111111010111", 410 => "01110001011101110111001101110111",411 => "01101110001010110010111000101011", 412 => "01011101000000000101111100000000", 413 => "01110111101111010111010110111101", 414 => "00010111010110111001011101011011", 415 => "01101011111010010110101111101000", 416 => "01010101011000100101010101110010"
																	,417 => "10111101100000001011110110010000", 418 => "01011100100111000101110010001100", 419 => "01001011100111110100101110011010", 420 => "11011101111010011101110111101011", 421 => "11111110100000111101111000000011", 422 => "00111011100011110011101010000111", 423 => "00101110011110010010111001111001", 424 => "00010111101110000001011010111000", 425 => "00001011100111010000101110011100", 426 => "01011010111001100101101010101110", 427 => "10111011110101011011001111010101"
																	,428 => "10111110101001111011111010110111", 429 =>"01101101110011110110110111001011", 430 => "11111101111011000111110111101110", 431 => "00010101110001010001010111000100", 432 => "10101011110100011011101110010001", 433 => "00100101110000110010010101000111", 434 => "11011010111000011101101011100001", 435 => "01010101110100110101010101010011", 436 => "11101011100101000110101110010100", 437 => "00110101110101010011010111110001", 438 => "01010111001100110101001100110011", 439 => "11011101101010110101110110101011"
																	,440 => "10111110000000011011111000001001", 441 => "00101011101111000010101110110100", 442 => "10010111000011001001011100001001", 443 => "11011111101011011101111110101111", 444 => "11100101111110001100010101111000", 445 => "01100101110101000110010011011100", 446 => "00010111001001010001011100100101", 447 => "10001011101100011000101010110001", 448 => "10001011100010111000101110001010", 449 => "11101011101000011110101111101001", 450 => "11000001011100001100100101110000", 451 => "01011100100111010101110010011100"
																	,452 => "10111000001000011011100000110001", 453 => "10100101110110011010010111010001", 454 => "10010111011100101001011101110111", 455 => "11011110111011111101111011101101", 456 =>"01101110101111110111111011111111", 457 => "10011100101110111001110000111111", 458 =>"11111010111010111111101011101011", 459 =>"11101111011111011110111101011101", 460 =>"00010111001010110000011100101011", 461 => "11001010101110100100101010111110", 462 => "01111111011110100111111111111010", 463 =>"00101110100111100010011010011110", 464 =>"01000111101110110100011111111011", 465 => "01011111010100100101111101010000"
																	,466 => "10111011100000011011101110010001", 467 => "10100101110110011010010111010001", 468 => "01110111110110000111011111011101", 469 => "01010101110011010101010111001111", 470 =>"00100110101011000011011011101100", 471 => "11001010111010011100101001101101", 472 =>"00101110111010100010111011101010", 473 => "11110101110000011111010110000001", 474 => "11101110111100001010111011110000", 475 => "00101110010010100010111001011000", 476 => "10101111101110001010110110111000", 477 =>"10101110110100111000111011010011", 478 =>"01111011101110100111101010111010"
																	,479 =>"10111100010000101011110001000110", 480 => "11001110111101101100111011110010", 481 =>"11000101110010011000010111001000", 482 =>"00111011111101010111101111110101", 483 =>"00001111011111000000110101110100", 484 => "01010101110110001101010111001000", 485 => "00100111101111110010011110111111", 486 => "11011010111011101101101011111110", 487 => "11010111001110001100011100111000", 488 => "01001011110011110100101111001011", 489 => "01110111001000010111011110100001", 490 => "01011110110100110100111011010011", 491 => "01110111010101110111011001010111", 492 => "10000101111110111010010111111011", 493 => "10100101110100101110010111010010", 494 => "10001011100100011100101110010001", 495 => "11111010101101011111101011110101", 496 => "00100101111110110010010110111011"
																	,497 => "10111110110001011011111011010101", 498 => "10111011001111001011101100110100", 499 => "10111001100101101011100110010011",																	
																	500 => "00111110001001110011111000101111", 501 => "01110100111110010111010011110001", 502 => "11100010011101011110001001110111", 503 => "10011001111010001001100111101001", 504 => "10000101011111001001010100111100", 505 =>"11100111110011101110011011001100", 506 => "00111011101110000011101110111000", 507 => "00111000101101000011100011110100", 508 => "00111000101101110111100010110111", 509 => "11001111110001101100111011000111", 510 => "01001111100001110100101110000111", 511 => "01000011101010110000001110101011", 512 => "00100011100000000010101110000000", 513 => "01110001111011010011000111101101", 514 => "00001110010110111000111001011011", 515 => "01001111011010100100111101101000", 516 => "01010100010100100101010001110010"
																	,517 => "00111011000000000011101100100000", 518 => "00010001110111000001000111001100", 519 => "01000111000111110100011100011010", 520 => "11011100111010011101110011101011", 521 => "11100000011000111100000011100011", 522 => "00001111100011110000101110000111", 523 => "00111000011110010011100001111001", 524 => "00111000101110000011100110111000", 525 => "00111000000111010011100000011100", 526 => "00011110110010100001101011001110", 527 => "10011101110101011000110111010101"
																	,528 => "00111110100101110011111010110111", 529 =>"01100011110011110110001111001011", 530 => "11111001111011000111100111101110", 531 => "00010011100001010001001110000100", 532 => "01100010010111010111001000011101", 533 => "00011101000000110001111100000111", 534 => "00111110110000010011111011000001", 535 => "00011110100100110001111000010011", 536 => "00111111000101001011111100010100", 537 => "00011101100100110001111110010001", 538 => "01001110001100110100011000110011", 539 => "10100111101010111110011110101011"
																	,540 => "00111100000010010011111000001001", 541 => "00100110011111000010011001110100", 542 => "10000001110011001000000111001001", 543 => "11110001111011011111000111101111", 544 => "11100101100011101100010100001110", 545 => "00011111000101000001101100011100", 546 => "00111000001001010011100000100101", 547 => "00111100001100010011110100110001", 548 => "00111100000010110011110000001010", 549 => "00111111001011010011101100101001", 550 => "11001110000000001101111000000000", 551 => "00000111100111001000011110011100"
																	,552 => "00101000001100010011100000110001", 553 => "10100000111110011010000011110001", 554 => "10000011111100101000001111110111", 555 => "11000111111011111100011111101101", 556 =>"01101110001111110111111001111111", 557 => "10011100111000011001111011100101", 558 =>"00111111110010110011111111001011", 559 =>"11001111011111011100111101011101", 560 =>"00111000001010110010100000101011", 561 => "11001110010100101000111000010010", 562 => "00111011111110100011101011111010", 563 =>"00000111100111100000001110011110", 564 =>"01000011101110110100001010111011", 565 => "01100011110100000111001111010000"
																	,566 => "00101011100100010011101110010001", 567 => "10101001101111111010100110011111", 568 => "01110011110110000111001111011101", 569 => "01010001110011010101000111001111", 570 =>"00100100001111000011010001111100", 571 => "11001110010010011100110001001101", 572 =>"00111000111010100011100011101010", 573 => "00111111100000010011111111000001", 574 => "00111111011100000111111101110000", 575 => "00111000010010010011100101001000", 576 => "10011101101110001001100110111000", 577 =>"10011010001110111000101000111011", 578 =>"01001111110110100100101111011010"
																	,579 =>"00110100010001100011110001000110", 580 => "11001100111100111100110011110010", 581 =>"11000000111010011000000011101000", 582 =>"00111110001111010111111000111101", 583 =>"00001110100011110000110010000111", 584 => "01010011100110001101001111011000", 585 => "00111001001111110011100100111111", 586 => "10011110110011101001111011011110", 587 => "00111110001110000010111000111000", 588 => "00111010010011110111101000001111", 589 => "00111011001000010011101000100001", 590 => "00011110110100110001011011010011", 591 => "01100111010101110110001101010111", 592 => "10000001111110111001000111111011", 593 => "10100001110100101110000111010010", 594 => "10000111000100011001011100010001", 595 => "11111000111101011101100011110101", 596 => "00100111001110110010010100111011"
																	,597 => "00101110110101010011111011010101", 598 => "01100100111101010110010011110100", 599 => "00110010011110100011001001111111",																	
														      	600 => "01010110001011110101111000101111", 601 => "01011011101100011101101110110001", 602 => "01011111000101011101111100010111", 603 => "01011100111010000101110011101001", 604 => "01001100111011000101110010101100", 605 =>"01011111110011100101111011001100", 606 => "01011011101110000101101110111000", 607 => "01011000101101000101100010010100", 608 => "01011000101101110101101010110111", 609 => "01011111110001100101101111000111", 610 => "01011011100001110101100110000111",611 => "01011010001010110100101000101011", 612 => "01011001000000000101110100000000", 613 => "01011011101011010001101110101101", 614 => "01011000010110111101100001011011", 615 => "01011011011010100101101101101000", 616 => "01011010101000100001101010100010"
																	,617 => "01001011001000000101101100100000", 618 => "01011000100011001101100010001100", 619 => "01011010000111110101101000011010", 620 => "01011110111010010101111011101011", 621 => "01111110100000110101111000000011", 622 => "01011001100011110101110110000111", 623 => "01011000011110010101100001111001", 624 => "01011000101110000101100000111000", 625 => "01011000000111000101000000011100", 626 => "01011010110010100100101011001110", 627 => "01011101110101010101010111010101"
																	,628 => "01001110101101110101111010110111", 629 =>"01011011010010110111101101001011", 630 => "01011111111011001101111111101110", 631 => "01011000100001010101100010000100", 632 => "01001011110100010101101110010001", 633 => "01011001000000110101101100000111", 634 => "01011110110000010101111011000001", 635 => "01001011100100110100101111010011", 636 => "01011111000101000101101100010100", 637 => "01011001100100110101000110010001", 638 => "01011010001100110101111000110011", 639 => "01011101101010110111110110101011"
																	,640 => "01001110000010010101111000001001", 641 => "01011001001101001101100100110100", 642 => "01011100000011000101110000001001", 643 => "01011111101011010101111110101111", 644 => "01111110101010000101111000101000", 645 => "01011011000101000101111100011100", 646 => "01011000001001010101100000100101", 647 => "10010110001100011001011010110001", 648 => "01011100000010100101010000001010", 649 => "01011111001011010100111100101001", 650 => "01011110000000000101011000000000", 651 => "01011000100111000101100010011100"
																	,652 => "00000010001111110000011000111111", 653 => "01011101000100011101110100010001", 654 => "01011100011100110101110001110111", 655 => "01011110111011110101111011101101", 656 =>"01001011101111110101101111111111", 657 => "01011100111000010101111011100101", 658 =>"01011111110010110101111111001011", 659 =>"01011111011111010101111101101101", 660 =>"01011000001010110101100010101011", 661 => "01011110010100100101111101010010", 662 => "01011011111110100101101101111010", 663 =>"01011000100111100101101010011110", 664 =>"01011010001110110101101100111011", 665 => "01011011010100000101001101010000"
																	,666 => "01010011100100010101101110010001", 667 => "01011101010011111101110101001111", 668 => "01011011110110000101101111011101", 669 => "01011010100011010101101010001111", 670 =>"01001001111011000101100110101100", 671 => "01011110010010010101110001001101", 672 =>"01011000111010100101100011101010", 673 => "01011111100000010101111110100001", 674 => "01011111011100000101110101110000", 675 => "01011000010010010101110001001000", 676 => "01011101101110000101111110111000", 677 =>"01011100110100110101010011010011", 678 =>"01011011110110100101111111011010"
																	,679 =>"01011000010001100101110001000110", 680 => "01011110011100110101111001110010", 681 =>"10101110000010011110111000001000", 682 =>"01011001111101010001100111110101", 683 =>"01011010011011000101100001100100", 684 => "01011010100110001101101011011000", 685 => "01011001001111110101100100111111", 686 => "01011110110011100101111011000110", 687 => "01011110001110000101111010111000", 688 => "01011010010011110001101101001111", 689 => "01011011001000010101101110100001", 690 => "01011010110100110101111011010011", 691 => "01011011010101110101111101010111", 692 => "01011100001110110111110000111011", 693 => "01011101000100100111110100010010", 694 => "01011100010100010101110000010001", 695 => "01011111110101010101110111010101", 696 => "01011001001110110101100110111011"
																	,697 => "01010110110101010101111011010101", 698 => "01011011001101100101101100110100", 699 => "01011001100101100101100110010011",																	
												    				700 => "10010010001011111001011000101111", 701 => "10010011101100001001001110110001", 702 => "10010111000101010001011100010111", 703 => "10010100111010001001010011101001", 704 => "10000100111011001001010010101100", 705 =>"10010111110011101001010111001100", 706 => "10010011101110001001001110111000", 707 => "10010000101101001001000010010100", 708 => "10010000101101111001010010110111", 709 => "10010111110001111001001111000111", 710 => "10010011100001111001000110000111",711 => "10010010001010111001101000101011", 712 => "10010001000000001001100100000000", 713 => "10010011101011011101001110101101", 714 => "10010000010110111101000001011011", 715 => "10011011011010001001001101101000", 716 => "10010010101000001001001010100010"
																	,717 => "10000011001000001001001100100000", 718 => "10010000100001001001000010001100", 719 => "10010010000111111001001000011010", 720 => "10010110111010011001011011101011", 721 => "10110110100000111001011000000011", 722 => "10010001100011111001100110000111", 723 => "10010000011110011001000001111001", 724 => "10010000101110001001000000111000", 725 => "10010000000111001000000000011100", 726 => "10010010110011101000001011001110", 727 => "10010101110101011001110111010101"
																	,728 => "10000110101101111001011010110111", 729 =>"10010011010011111001001101001011", 730 => "10010111111011000001011111101110", 731 => "10010000100001011001000010000100", 732 => "10000011110100011001001110010001", 733 => "10010001000000111001010100000111", 734 => "10010110110000011001011011000001", 735 => "10010010100100111001001011010011", 736 => "10010111000101001001111100010100", 737 => "10010001100100011001100110010001", 738 => "10010010001100111001011000110011", 739 => "10010101101010111000010110101011"
																	,740 => "10000110000010011001011000001001", 741 => "10010001001111001001000100110100", 742 => "10010100000011001001010000001001", 743 => "10010111101011011001011110101111", 744 => "10110110101010001001011000101000", 745 => "10010011000101001001101100011100", 746 => "10010000001001011001000000100101", 747 => "10010100001100011001010010110001", 748 => "10010100000010101100010000001010", 749 => "10010111001010011000011100101001", 750 => "10010110000000001001111000000000", 751 => "10010000100111001011000010011100"
																	,752 => "10000000001100011001000000110001", 753 => "10010101001100011001010100010001", 754 => "10010100011100101001010001110111", 755 => "10010110111011111001011011101101", 756 =>"10000011101111111001001111111111", 757 => "10010100111000011001000011100101", 758 =>"10010111110010111001011111001011", 759 =>"10010111011111011001011101101101", 760 =>"10010000001010111001010000101011", 761 => "10010110010100101001011101010010", 762 => "10010011111110101001001101111010", 763 =>"10010000100111101001000110011110", 764 =>"10010010001110111001011000111011", 765 => "10010011010100001101001101010000"
																	,766 => "10000011100100011001001110010001", 767 => "10010101010111111001010101001111", 768 => "10010011110110001001001111011101", 769 => "10010010100011011001001010001111", 770 =>"10000001111011001001000110101100", 771 => "10010110010010011001001001001101", 772 =>"10010000111010101001000011101010", 773 => "10010111100000011001011110100001", 774 => "10010111011100001000011101110000", 775 => "10010000010010001001010001001000", 776 => "10010101101110001001011110111000", 777 =>"10010100110100111001000011010011", 778 =>"10010011110110101000001111011010"
																	,779 =>"10010100010001101001010001000110", 780 => "10010110011101101001011001110010", 781 =>"10010110000010011101011000001000", 782 =>"10010001111101011101000111110101", 783 =>"10010010011011001001000001100100", 784 => "10010010100110000001001000011000", 785 => "10010001001111111001000100111111", 786 => "10010110110011101001011011000110", 787 => "10010110001110001001001000111000", 788 => "10010010010011111001001101001111", 789 => "10010011001000011001001110100001", 790 => "10010010110100111001000011010011", 791 => "01101001101010111101001101010111", 792 => "10010100001110111101010000111011", 793 => "10010101000100101011010100010010", 794 => "10010100100100011001010000010001", 795 => "10010111110101011001011011010101", 796 => "10010001001110111001010100111011"
																	,797 => "10000110110101011001011011010101", 798 => "10010011001111001001001100110100", 799 => "10010001100101101001000110010011",																
																	800 => "10000110001011111001011000101111", 801 => "10010011101110011001001110110001", 802 => "11001011000101010100101100010111", 803 => "10010100111010001001010011101001", 804 => "10000100111011001001010010101100", 805 =>"10010111010011001001010111001100", 806 => "10010011101110001001001110111000", 807 => "10010000101101001001000010110000", 808 => "10010000101101111001010010110111", 809 => "10010111110001111001001111000111", 810 => "10010011100001111001000110000111",811 => "10010010001010111001000000101011", 812 => "10010001000000001001010100000000", 813 => "10010011101111011001001110101101", 814 => "10010000010110111101000001011011", 815 => "10010011011010101001001101101000", 816 => "10010010101000101001101010100010"
																	,817 => "10000011001000001001001100100000", 818 => "10010000100111001001000010001100", 819 => "10010010000111111001001000011010", 820 => "10010110111010011001011011101011", 821 => "10110110100000111001011000000011", 822 => "10010011100001111001100110000111", 823 => "10010000011110011001000001111001", 824 => "10010000101110001001000010101000", 825 => "10010000000111001000000000011100", 826 => "10010010110011101000001011001110", 827 => "10010101110101011001110111010101"
																	,828 => "10000110101101111001011010110111", 829 =>"10010011010011111001001101001011", 830 => "10010111111011000001011111101110", 831 => "10010000100001011001000010000100", 832 => "10000011110100011001001110010001", 833 => "10010000000001111001010100000111", 834 => "10010110110000011001011011000001", 835 => "10010010100100111001001010011011", 836 => "10010111000101001001111100010100", 837 => "10010001100100011001100110010001", 838 => "10010010001100111001110001100110", 839 => "10010101101010111001110110101011"
																	,840 => "10000110000010011001011000001001", 841 => "10010001001111001001000100110100", 842 => "10010100000011001001010000001001", 843 => "10010111101011011001011110101111", 844 => "10110110101010001001011000101000", 845 => "10010001000111001001101100011100", 846 => "10010000001001011001000000100101", 847 => "10010100001100011001010000100001", 848 => "10010100000010101000010000001010", 849 => "10010111001010011000011100101001", 850 => "10010110000000001000011000000000", 851 => "10010000100111001011000010011100"
																	,852 => "10000000001100011001000000110001", 853 => "10010101000110011001010100010001", 854 => "10010100011100101001010001110111", 855 => "10010110111011111001011011101101", 856 =>"10000011101111111001001111111111", 857 => "10010101111001011001000011100101", 858 =>"10010111110010111001011111001011", 859 =>"10010111011111011001011101111111", 860 =>"10010000001010111001000100101011", 861 => "10010110010100101001011101010010", 862 => "10010011111110101001001011111010", 863 =>"10010000100111101001000110011110", 864 =>"10010010001110111001001010111011", 865 => "10010011010101001001001101010000"
																	,866 => "10000011100100011001001110010001", 867 => "10010101010111111001010101001111", 868 => "10010011110110001001001111011101", 869 => "10010010100011011001001010001111", 870 =>"10000001111011001001000110101100", 871 => "10010111010011011001001001001101", 872 =>"10010000111010101001000011101010", 873 => "10010111100000011001011110000101", 874 => "10010111011100001001001101110000", 875 => "10010000010010001001010001001000", 876 => "10010101101110001001000110111000", 877 =>"10010100110100111001000011010011", 878 =>"10010011110110101001000111011010"
																	,879 =>"10000100010001101001010001000110", 880 => "10010110011101101001011001110010", 881 =>"10010110000010010001011000001000", 882 =>"10010001111101011101000111110101", 883 =>"10010010011011001001000001100100", 884 => "10010010101110001001001000011000", 885 => "10010001001111111001000100111111", 886 => "10010110110011101001011011001111", 887 => "10010110001110001001011100111000", 888 => "10010010010011111001001101001111", 889 => "10010011001000011001001000100001", 890 => "10010010110100111001000011010011", 891 => "10010011010101111001000101010111", 892 => "10010100001111111001010000111011", 893 => "10010101000100101011010100010010", 894 => "10010100000110011001010000010001", 895 => "10010111110101011001011011010101", 896 => "10010001001110111001010100111011"
																	,897 => "10000110110101011001011011010101", 898 => "10010011001111001001001100110100", 899 => "10010001100101101001000110010011",
																	900 => "00000110001011110000111000101111", 901 => "01110110001010010111011000100001", 902 => "11100010111000110110001011100001", 903 => "10011101001000001001110100100001", 904 => "10000111110000011001010110000001", 905 =>"00001111110011000000110111001100", 906 => "01110111000000010111011100000001", 907 => "00010110100000010001011010000101", 908 => "00001000101101110010100010110111", 909 => "11100001110001111110100111000111", 910 => "00001011100001110000111110000111",911 => "00001010001010110000111000101011", 912 => "00000101000000000000000100000000", 913 => "00001011101111010000101110101101", 914 => "00001000010110110010100001011011", 915 => "00001011011010001000101101101000", 916 => "00001010101000101000101010100010"
																	,917 => "00000011001000000000101100100000", 918 => "00010001100100010001000110000001", 919 => "11100010111001001110001011100001", 920 => "11011101011000111101110101100001", 921 => "11100100111000011100000001100001", 922 => "00001001100001110000000110000111", 923 => "00001111001000010000111100100001", 924 => "00010111000000010001011100010001", 925 => "00001000000111001000100000011100", 926 => "01000010110011100110001011001110", 927 => "10000101110101011001010111010101"
																	,928 => "00000110101101110000111010110111", 929 =>"01101001011010010110100101100001", 930 => "11111101110000110111110111000001", 931 => "00010000100000000001000010000001", 932 => "01100110011000010111001000100001", 933 => "00001001000001110000110100000111", 934 => "11011000001000011101100000100001", 935 => "01010010011000010101001001101001", 936 => "00001111000101000100111100010100", 937 => "00000101100100010001010110010001", 938 => "00001010001100110000001000110011", 939 => "00001101101010110001110110101011"
																	,940 => "00000110000010010000111000001001", 941 => "00100110100100010010011010000001", 942 => "10000001001001001000000100100001", 943 => "11110101111000111111010111100001", 944 => "11101101100000011100010100000001", 945 => "00001011000111000000001100011100", 946 => "00000100101000010000010010100001", 947 => "10000110001000011000011000110001", 948 => "00001100000010101000110000001010", 949 => "00001111001010010010111100101001", 950 => "00001110000000000001111000000000", 951 => "00001000100111000010100010011100"
																	,952 => "00000000001100010000100000110001", 953 => "10100010001100011010001000100001", 954 => "10001110111001001000111011100001", 955 => "11011101101000111101110110100001", 956 =>"01101011101000010111111111100001", 957 => "00001100111001010000100011100101", 958 =>"11111001011000011111100101100001", 959 =>"11101111101000011110111110100011", 960 =>"00001000001010110000000000101011", 961 => "00001110010100100000110001010010", 962 => "00001011111110100000101011111010", 963 =>"00001000100111100000100110011110", 964 =>"01000010001110110100001000011011", 965 => "10000101101010001000101101010000"
																	,966 => "00000011100100010000101110010001", 967 => "10101001111100011010100111100001", 968 => "01111011101001000111101110100001", 969 => "01010001111000110101000111100001", 970 =>"00100001110000010011010110000001", 971 => "00001110010011010000101001001101", 972 =>"00011101010000010001110101000001", 973 => "11110000001000011111000000100101", 974 => "00001111011100000010111101110000", 975 => "00001000010010000000000001001000", 976 => "00001101101110000000100110111000", 977 =>"00001100110100110000100011010011", 978 =>"00000111110110100000011101011010"
																	,979 =>"00001000010001100000110001000110", 980 => "11001110011000011100111001000001", 981 =>"11000001000000001000000100000001", 982 =>"00111110101000010111111010100001", 983 =>"00001110000010010000110010000001", 984 => "00001010100110000000101000011000", 985 => "00100111111000010010011111100001", 986 => "11011001110000011101100111000000", 987 => "00001110001110000000011000111000", 988 => "00001010010011110000100001001111", 989 => "00001011001000010000101000100001", 990 => "00001010110100110000100011010011", 991 => "00000111010101110000011111010111", 992 => "00001100001110110100110000111011", 993 => "00001101000100100010110100010010", 994 => "00001100100100010000110000010001", 995 => "00001111110101010000111011010101", 996 => "00001001001110110100100100111011"
																	,997 => "00000110110101010000111011010101", 998 => "01100110110000101100110100010011", 999 => "00110010011000100011001001100001");

begin

	process(clock)
	variable index_Input:integer;
	begin
		index_Input := 0;
		for i in 0 to 999 loop
			if(VAdress(i) = VirtualAddress) then
				index_Input:= i;
			end if; 
		end loop;
		PhysicalAddressOut<= PAdress(index_Input);
		if(cache_type = '0') then
			outputData(31 downto 0 )<=DataOutput1(index_Input);
			outputData(63 downto 32)<=DataOutput2(index_Input);
		else
			outputData(31 downto 0 )<=DataOutput1(index_Input);
			outputData(63 downto 32)<="UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU";
		end if;
	end process;
end Behavioral;

